magic
tech sky130A
magscale 1 2
timestamp 1635172635
<< obsli1 >>
rect 1104 2159 418876 417809
<< obsm1 >>
rect 382 2128 419506 417840
<< metal2 >>
rect 1858 419200 1914 420000
rect 5538 419200 5594 420000
rect 9218 419200 9274 420000
rect 12898 419200 12954 420000
rect 16578 419200 16634 420000
rect 20258 419200 20314 420000
rect 23938 419200 23994 420000
rect 27618 419200 27674 420000
rect 31298 419200 31354 420000
rect 34978 419200 35034 420000
rect 38658 419200 38714 420000
rect 42338 419200 42394 420000
rect 46018 419200 46074 420000
rect 49698 419200 49754 420000
rect 53378 419200 53434 420000
rect 57058 419200 57114 420000
rect 60738 419200 60794 420000
rect 64418 419200 64474 420000
rect 68098 419200 68154 420000
rect 71778 419200 71834 420000
rect 75458 419200 75514 420000
rect 79138 419200 79194 420000
rect 82818 419200 82874 420000
rect 86590 419200 86646 420000
rect 90270 419200 90326 420000
rect 93950 419200 94006 420000
rect 97630 419200 97686 420000
rect 101310 419200 101366 420000
rect 104990 419200 105046 420000
rect 108670 419200 108726 420000
rect 112350 419200 112406 420000
rect 116030 419200 116086 420000
rect 119710 419200 119766 420000
rect 123390 419200 123446 420000
rect 127070 419200 127126 420000
rect 130750 419200 130806 420000
rect 134430 419200 134486 420000
rect 138110 419200 138166 420000
rect 141790 419200 141846 420000
rect 145470 419200 145526 420000
rect 149150 419200 149206 420000
rect 152830 419200 152886 420000
rect 156510 419200 156566 420000
rect 160190 419200 160246 420000
rect 163870 419200 163926 420000
rect 167550 419200 167606 420000
rect 171322 419200 171378 420000
rect 175002 419200 175058 420000
rect 178682 419200 178738 420000
rect 182362 419200 182418 420000
rect 186042 419200 186098 420000
rect 189722 419200 189778 420000
rect 193402 419200 193458 420000
rect 197082 419200 197138 420000
rect 200762 419200 200818 420000
rect 204442 419200 204498 420000
rect 208122 419200 208178 420000
rect 211802 419200 211858 420000
rect 215482 419200 215538 420000
rect 219162 419200 219218 420000
rect 222842 419200 222898 420000
rect 226522 419200 226578 420000
rect 230202 419200 230258 420000
rect 233882 419200 233938 420000
rect 237562 419200 237618 420000
rect 241242 419200 241298 420000
rect 244922 419200 244978 420000
rect 248602 419200 248658 420000
rect 252282 419200 252338 420000
rect 256054 419200 256110 420000
rect 259734 419200 259790 420000
rect 263414 419200 263470 420000
rect 267094 419200 267150 420000
rect 270774 419200 270830 420000
rect 274454 419200 274510 420000
rect 278134 419200 278190 420000
rect 281814 419200 281870 420000
rect 285494 419200 285550 420000
rect 289174 419200 289230 420000
rect 292854 419200 292910 420000
rect 296534 419200 296590 420000
rect 300214 419200 300270 420000
rect 303894 419200 303950 420000
rect 307574 419200 307630 420000
rect 311254 419200 311310 420000
rect 314934 419200 314990 420000
rect 318614 419200 318670 420000
rect 322294 419200 322350 420000
rect 325974 419200 326030 420000
rect 329654 419200 329710 420000
rect 333334 419200 333390 420000
rect 337014 419200 337070 420000
rect 340786 419200 340842 420000
rect 344466 419200 344522 420000
rect 348146 419200 348202 420000
rect 351826 419200 351882 420000
rect 355506 419200 355562 420000
rect 359186 419200 359242 420000
rect 362866 419200 362922 420000
rect 366546 419200 366602 420000
rect 370226 419200 370282 420000
rect 373906 419200 373962 420000
rect 377586 419200 377642 420000
rect 381266 419200 381322 420000
rect 384946 419200 385002 420000
rect 388626 419200 388682 420000
rect 392306 419200 392362 420000
rect 395986 419200 396042 420000
rect 399666 419200 399722 420000
rect 403346 419200 403402 420000
rect 407026 419200 407082 420000
rect 410706 419200 410762 420000
rect 414386 419200 414442 420000
rect 418066 419200 418122 420000
rect 386 0 442 800
rect 1214 0 1270 800
rect 2042 0 2098 800
rect 2870 0 2926 800
rect 3790 0 3846 800
rect 4618 0 4674 800
rect 5446 0 5502 800
rect 6274 0 6330 800
rect 7194 0 7250 800
rect 8022 0 8078 800
rect 8850 0 8906 800
rect 9678 0 9734 800
rect 10598 0 10654 800
rect 11426 0 11482 800
rect 12254 0 12310 800
rect 13082 0 13138 800
rect 14002 0 14058 800
rect 14830 0 14886 800
rect 15658 0 15714 800
rect 16486 0 16542 800
rect 17406 0 17462 800
rect 18234 0 18290 800
rect 19062 0 19118 800
rect 19890 0 19946 800
rect 20810 0 20866 800
rect 21638 0 21694 800
rect 22466 0 22522 800
rect 23386 0 23442 800
rect 24214 0 24270 800
rect 25042 0 25098 800
rect 25870 0 25926 800
rect 26790 0 26846 800
rect 27618 0 27674 800
rect 28446 0 28502 800
rect 29274 0 29330 800
rect 30194 0 30250 800
rect 31022 0 31078 800
rect 31850 0 31906 800
rect 32678 0 32734 800
rect 33598 0 33654 800
rect 34426 0 34482 800
rect 35254 0 35310 800
rect 36082 0 36138 800
rect 37002 0 37058 800
rect 37830 0 37886 800
rect 38658 0 38714 800
rect 39486 0 39542 800
rect 40406 0 40462 800
rect 41234 0 41290 800
rect 42062 0 42118 800
rect 42890 0 42946 800
rect 43810 0 43866 800
rect 44638 0 44694 800
rect 45466 0 45522 800
rect 46386 0 46442 800
rect 47214 0 47270 800
rect 48042 0 48098 800
rect 48870 0 48926 800
rect 49790 0 49846 800
rect 50618 0 50674 800
rect 51446 0 51502 800
rect 52274 0 52330 800
rect 53194 0 53250 800
rect 54022 0 54078 800
rect 54850 0 54906 800
rect 55678 0 55734 800
rect 56598 0 56654 800
rect 57426 0 57482 800
rect 58254 0 58310 800
rect 59082 0 59138 800
rect 60002 0 60058 800
rect 60830 0 60886 800
rect 61658 0 61714 800
rect 62486 0 62542 800
rect 63406 0 63462 800
rect 64234 0 64290 800
rect 65062 0 65118 800
rect 65890 0 65946 800
rect 66810 0 66866 800
rect 67638 0 67694 800
rect 68466 0 68522 800
rect 69386 0 69442 800
rect 70214 0 70270 800
rect 71042 0 71098 800
rect 71870 0 71926 800
rect 72790 0 72846 800
rect 73618 0 73674 800
rect 74446 0 74502 800
rect 75274 0 75330 800
rect 76194 0 76250 800
rect 77022 0 77078 800
rect 77850 0 77906 800
rect 78678 0 78734 800
rect 79598 0 79654 800
rect 80426 0 80482 800
rect 81254 0 81310 800
rect 82082 0 82138 800
rect 83002 0 83058 800
rect 83830 0 83886 800
rect 84658 0 84714 800
rect 85486 0 85542 800
rect 86406 0 86462 800
rect 87234 0 87290 800
rect 88062 0 88118 800
rect 88982 0 89038 800
rect 89810 0 89866 800
rect 90638 0 90694 800
rect 91466 0 91522 800
rect 92386 0 92442 800
rect 93214 0 93270 800
rect 94042 0 94098 800
rect 94870 0 94926 800
rect 95790 0 95846 800
rect 96618 0 96674 800
rect 97446 0 97502 800
rect 98274 0 98330 800
rect 99194 0 99250 800
rect 100022 0 100078 800
rect 100850 0 100906 800
rect 101678 0 101734 800
rect 102598 0 102654 800
rect 103426 0 103482 800
rect 104254 0 104310 800
rect 105082 0 105138 800
rect 106002 0 106058 800
rect 106830 0 106886 800
rect 107658 0 107714 800
rect 108486 0 108542 800
rect 109406 0 109462 800
rect 110234 0 110290 800
rect 111062 0 111118 800
rect 111982 0 112038 800
rect 112810 0 112866 800
rect 113638 0 113694 800
rect 114466 0 114522 800
rect 115386 0 115442 800
rect 116214 0 116270 800
rect 117042 0 117098 800
rect 117870 0 117926 800
rect 118790 0 118846 800
rect 119618 0 119674 800
rect 120446 0 120502 800
rect 121274 0 121330 800
rect 122194 0 122250 800
rect 123022 0 123078 800
rect 123850 0 123906 800
rect 124678 0 124734 800
rect 125598 0 125654 800
rect 126426 0 126482 800
rect 127254 0 127310 800
rect 128082 0 128138 800
rect 129002 0 129058 800
rect 129830 0 129886 800
rect 130658 0 130714 800
rect 131486 0 131542 800
rect 132406 0 132462 800
rect 133234 0 133290 800
rect 134062 0 134118 800
rect 134982 0 135038 800
rect 135810 0 135866 800
rect 136638 0 136694 800
rect 137466 0 137522 800
rect 138386 0 138442 800
rect 139214 0 139270 800
rect 140042 0 140098 800
rect 140870 0 140926 800
rect 141790 0 141846 800
rect 142618 0 142674 800
rect 143446 0 143502 800
rect 144274 0 144330 800
rect 145194 0 145250 800
rect 146022 0 146078 800
rect 146850 0 146906 800
rect 147678 0 147734 800
rect 148598 0 148654 800
rect 149426 0 149482 800
rect 150254 0 150310 800
rect 151082 0 151138 800
rect 152002 0 152058 800
rect 152830 0 152886 800
rect 153658 0 153714 800
rect 154486 0 154542 800
rect 155406 0 155462 800
rect 156234 0 156290 800
rect 157062 0 157118 800
rect 157982 0 158038 800
rect 158810 0 158866 800
rect 159638 0 159694 800
rect 160466 0 160522 800
rect 161386 0 161442 800
rect 162214 0 162270 800
rect 163042 0 163098 800
rect 163870 0 163926 800
rect 164790 0 164846 800
rect 165618 0 165674 800
rect 166446 0 166502 800
rect 167274 0 167330 800
rect 168194 0 168250 800
rect 169022 0 169078 800
rect 169850 0 169906 800
rect 170678 0 170734 800
rect 171598 0 171654 800
rect 172426 0 172482 800
rect 173254 0 173310 800
rect 174082 0 174138 800
rect 175002 0 175058 800
rect 175830 0 175886 800
rect 176658 0 176714 800
rect 177578 0 177634 800
rect 178406 0 178462 800
rect 179234 0 179290 800
rect 180062 0 180118 800
rect 180982 0 181038 800
rect 181810 0 181866 800
rect 182638 0 182694 800
rect 183466 0 183522 800
rect 184386 0 184442 800
rect 185214 0 185270 800
rect 186042 0 186098 800
rect 186870 0 186926 800
rect 187790 0 187846 800
rect 188618 0 188674 800
rect 189446 0 189502 800
rect 190274 0 190330 800
rect 191194 0 191250 800
rect 192022 0 192078 800
rect 192850 0 192906 800
rect 193678 0 193734 800
rect 194598 0 194654 800
rect 195426 0 195482 800
rect 196254 0 196310 800
rect 197082 0 197138 800
rect 198002 0 198058 800
rect 198830 0 198886 800
rect 199658 0 199714 800
rect 200578 0 200634 800
rect 201406 0 201462 800
rect 202234 0 202290 800
rect 203062 0 203118 800
rect 203982 0 204038 800
rect 204810 0 204866 800
rect 205638 0 205694 800
rect 206466 0 206522 800
rect 207386 0 207442 800
rect 208214 0 208270 800
rect 209042 0 209098 800
rect 209870 0 209926 800
rect 210790 0 210846 800
rect 211618 0 211674 800
rect 212446 0 212502 800
rect 213274 0 213330 800
rect 214194 0 214250 800
rect 215022 0 215078 800
rect 215850 0 215906 800
rect 216678 0 216734 800
rect 217598 0 217654 800
rect 218426 0 218482 800
rect 219254 0 219310 800
rect 220082 0 220138 800
rect 221002 0 221058 800
rect 221830 0 221886 800
rect 222658 0 222714 800
rect 223578 0 223634 800
rect 224406 0 224462 800
rect 225234 0 225290 800
rect 226062 0 226118 800
rect 226982 0 227038 800
rect 227810 0 227866 800
rect 228638 0 228694 800
rect 229466 0 229522 800
rect 230386 0 230442 800
rect 231214 0 231270 800
rect 232042 0 232098 800
rect 232870 0 232926 800
rect 233790 0 233846 800
rect 234618 0 234674 800
rect 235446 0 235502 800
rect 236274 0 236330 800
rect 237194 0 237250 800
rect 238022 0 238078 800
rect 238850 0 238906 800
rect 239678 0 239734 800
rect 240598 0 240654 800
rect 241426 0 241482 800
rect 242254 0 242310 800
rect 243082 0 243138 800
rect 244002 0 244058 800
rect 244830 0 244886 800
rect 245658 0 245714 800
rect 246578 0 246634 800
rect 247406 0 247462 800
rect 248234 0 248290 800
rect 249062 0 249118 800
rect 249982 0 250038 800
rect 250810 0 250866 800
rect 251638 0 251694 800
rect 252466 0 252522 800
rect 253386 0 253442 800
rect 254214 0 254270 800
rect 255042 0 255098 800
rect 255870 0 255926 800
rect 256790 0 256846 800
rect 257618 0 257674 800
rect 258446 0 258502 800
rect 259274 0 259330 800
rect 260194 0 260250 800
rect 261022 0 261078 800
rect 261850 0 261906 800
rect 262678 0 262734 800
rect 263598 0 263654 800
rect 264426 0 264482 800
rect 265254 0 265310 800
rect 266174 0 266230 800
rect 267002 0 267058 800
rect 267830 0 267886 800
rect 268658 0 268714 800
rect 269578 0 269634 800
rect 270406 0 270462 800
rect 271234 0 271290 800
rect 272062 0 272118 800
rect 272982 0 273038 800
rect 273810 0 273866 800
rect 274638 0 274694 800
rect 275466 0 275522 800
rect 276386 0 276442 800
rect 277214 0 277270 800
rect 278042 0 278098 800
rect 278870 0 278926 800
rect 279790 0 279846 800
rect 280618 0 280674 800
rect 281446 0 281502 800
rect 282274 0 282330 800
rect 283194 0 283250 800
rect 284022 0 284078 800
rect 284850 0 284906 800
rect 285678 0 285734 800
rect 286598 0 286654 800
rect 287426 0 287482 800
rect 288254 0 288310 800
rect 289174 0 289230 800
rect 290002 0 290058 800
rect 290830 0 290886 800
rect 291658 0 291714 800
rect 292578 0 292634 800
rect 293406 0 293462 800
rect 294234 0 294290 800
rect 295062 0 295118 800
rect 295982 0 296038 800
rect 296810 0 296866 800
rect 297638 0 297694 800
rect 298466 0 298522 800
rect 299386 0 299442 800
rect 300214 0 300270 800
rect 301042 0 301098 800
rect 301870 0 301926 800
rect 302790 0 302846 800
rect 303618 0 303674 800
rect 304446 0 304502 800
rect 305274 0 305330 800
rect 306194 0 306250 800
rect 307022 0 307078 800
rect 307850 0 307906 800
rect 308678 0 308734 800
rect 309598 0 309654 800
rect 310426 0 310482 800
rect 311254 0 311310 800
rect 312174 0 312230 800
rect 313002 0 313058 800
rect 313830 0 313886 800
rect 314658 0 314714 800
rect 315578 0 315634 800
rect 316406 0 316462 800
rect 317234 0 317290 800
rect 318062 0 318118 800
rect 318982 0 319038 800
rect 319810 0 319866 800
rect 320638 0 320694 800
rect 321466 0 321522 800
rect 322386 0 322442 800
rect 323214 0 323270 800
rect 324042 0 324098 800
rect 324870 0 324926 800
rect 325790 0 325846 800
rect 326618 0 326674 800
rect 327446 0 327502 800
rect 328274 0 328330 800
rect 329194 0 329250 800
rect 330022 0 330078 800
rect 330850 0 330906 800
rect 331678 0 331734 800
rect 332598 0 332654 800
rect 333426 0 333482 800
rect 334254 0 334310 800
rect 335174 0 335230 800
rect 336002 0 336058 800
rect 336830 0 336886 800
rect 337658 0 337714 800
rect 338578 0 338634 800
rect 339406 0 339462 800
rect 340234 0 340290 800
rect 341062 0 341118 800
rect 341982 0 342038 800
rect 342810 0 342866 800
rect 343638 0 343694 800
rect 344466 0 344522 800
rect 345386 0 345442 800
rect 346214 0 346270 800
rect 347042 0 347098 800
rect 347870 0 347926 800
rect 348790 0 348846 800
rect 349618 0 349674 800
rect 350446 0 350502 800
rect 351274 0 351330 800
rect 352194 0 352250 800
rect 353022 0 353078 800
rect 353850 0 353906 800
rect 354770 0 354826 800
rect 355598 0 355654 800
rect 356426 0 356482 800
rect 357254 0 357310 800
rect 358174 0 358230 800
rect 359002 0 359058 800
rect 359830 0 359886 800
rect 360658 0 360714 800
rect 361578 0 361634 800
rect 362406 0 362462 800
rect 363234 0 363290 800
rect 364062 0 364118 800
rect 364982 0 365038 800
rect 365810 0 365866 800
rect 366638 0 366694 800
rect 367466 0 367522 800
rect 368386 0 368442 800
rect 369214 0 369270 800
rect 370042 0 370098 800
rect 370870 0 370926 800
rect 371790 0 371846 800
rect 372618 0 372674 800
rect 373446 0 373502 800
rect 374274 0 374330 800
rect 375194 0 375250 800
rect 376022 0 376078 800
rect 376850 0 376906 800
rect 377770 0 377826 800
rect 378598 0 378654 800
rect 379426 0 379482 800
rect 380254 0 380310 800
rect 381174 0 381230 800
rect 382002 0 382058 800
rect 382830 0 382886 800
rect 383658 0 383714 800
rect 384578 0 384634 800
rect 385406 0 385462 800
rect 386234 0 386290 800
rect 387062 0 387118 800
rect 387982 0 388038 800
rect 388810 0 388866 800
rect 389638 0 389694 800
rect 390466 0 390522 800
rect 391386 0 391442 800
rect 392214 0 392270 800
rect 393042 0 393098 800
rect 393870 0 393926 800
rect 394790 0 394846 800
rect 395618 0 395674 800
rect 396446 0 396502 800
rect 397274 0 397330 800
rect 398194 0 398250 800
rect 399022 0 399078 800
rect 399850 0 399906 800
rect 400770 0 400826 800
rect 401598 0 401654 800
rect 402426 0 402482 800
rect 403254 0 403310 800
rect 404174 0 404230 800
rect 405002 0 405058 800
rect 405830 0 405886 800
rect 406658 0 406714 800
rect 407578 0 407634 800
rect 408406 0 408462 800
rect 409234 0 409290 800
rect 410062 0 410118 800
rect 410982 0 411038 800
rect 411810 0 411866 800
rect 412638 0 412694 800
rect 413466 0 413522 800
rect 414386 0 414442 800
rect 415214 0 415270 800
rect 416042 0 416098 800
rect 416870 0 416926 800
rect 417790 0 417846 800
rect 418618 0 418674 800
rect 419446 0 419502 800
<< obsm2 >>
rect 388 419144 1802 419200
rect 1970 419144 5482 419200
rect 5650 419144 9162 419200
rect 9330 419144 12842 419200
rect 13010 419144 16522 419200
rect 16690 419144 20202 419200
rect 20370 419144 23882 419200
rect 24050 419144 27562 419200
rect 27730 419144 31242 419200
rect 31410 419144 34922 419200
rect 35090 419144 38602 419200
rect 38770 419144 42282 419200
rect 42450 419144 45962 419200
rect 46130 419144 49642 419200
rect 49810 419144 53322 419200
rect 53490 419144 57002 419200
rect 57170 419144 60682 419200
rect 60850 419144 64362 419200
rect 64530 419144 68042 419200
rect 68210 419144 71722 419200
rect 71890 419144 75402 419200
rect 75570 419144 79082 419200
rect 79250 419144 82762 419200
rect 82930 419144 86534 419200
rect 86702 419144 90214 419200
rect 90382 419144 93894 419200
rect 94062 419144 97574 419200
rect 97742 419144 101254 419200
rect 101422 419144 104934 419200
rect 105102 419144 108614 419200
rect 108782 419144 112294 419200
rect 112462 419144 115974 419200
rect 116142 419144 119654 419200
rect 119822 419144 123334 419200
rect 123502 419144 127014 419200
rect 127182 419144 130694 419200
rect 130862 419144 134374 419200
rect 134542 419144 138054 419200
rect 138222 419144 141734 419200
rect 141902 419144 145414 419200
rect 145582 419144 149094 419200
rect 149262 419144 152774 419200
rect 152942 419144 156454 419200
rect 156622 419144 160134 419200
rect 160302 419144 163814 419200
rect 163982 419144 167494 419200
rect 167662 419144 171266 419200
rect 171434 419144 174946 419200
rect 175114 419144 178626 419200
rect 178794 419144 182306 419200
rect 182474 419144 185986 419200
rect 186154 419144 189666 419200
rect 189834 419144 193346 419200
rect 193514 419144 197026 419200
rect 197194 419144 200706 419200
rect 200874 419144 204386 419200
rect 204554 419144 208066 419200
rect 208234 419144 211746 419200
rect 211914 419144 215426 419200
rect 215594 419144 219106 419200
rect 219274 419144 222786 419200
rect 222954 419144 226466 419200
rect 226634 419144 230146 419200
rect 230314 419144 233826 419200
rect 233994 419144 237506 419200
rect 237674 419144 241186 419200
rect 241354 419144 244866 419200
rect 245034 419144 248546 419200
rect 248714 419144 252226 419200
rect 252394 419144 255998 419200
rect 256166 419144 259678 419200
rect 259846 419144 263358 419200
rect 263526 419144 267038 419200
rect 267206 419144 270718 419200
rect 270886 419144 274398 419200
rect 274566 419144 278078 419200
rect 278246 419144 281758 419200
rect 281926 419144 285438 419200
rect 285606 419144 289118 419200
rect 289286 419144 292798 419200
rect 292966 419144 296478 419200
rect 296646 419144 300158 419200
rect 300326 419144 303838 419200
rect 304006 419144 307518 419200
rect 307686 419144 311198 419200
rect 311366 419144 314878 419200
rect 315046 419144 318558 419200
rect 318726 419144 322238 419200
rect 322406 419144 325918 419200
rect 326086 419144 329598 419200
rect 329766 419144 333278 419200
rect 333446 419144 336958 419200
rect 337126 419144 340730 419200
rect 340898 419144 344410 419200
rect 344578 419144 348090 419200
rect 348258 419144 351770 419200
rect 351938 419144 355450 419200
rect 355618 419144 359130 419200
rect 359298 419144 362810 419200
rect 362978 419144 366490 419200
rect 366658 419144 370170 419200
rect 370338 419144 373850 419200
rect 374018 419144 377530 419200
rect 377698 419144 381210 419200
rect 381378 419144 384890 419200
rect 385058 419144 388570 419200
rect 388738 419144 392250 419200
rect 392418 419144 395930 419200
rect 396098 419144 399610 419200
rect 399778 419144 403290 419200
rect 403458 419144 406970 419200
rect 407138 419144 410650 419200
rect 410818 419144 414330 419200
rect 414498 419144 418010 419200
rect 418178 419144 419500 419200
rect 388 856 419500 419144
rect 498 734 1158 856
rect 1326 734 1986 856
rect 2154 734 2814 856
rect 2982 734 3734 856
rect 3902 734 4562 856
rect 4730 734 5390 856
rect 5558 734 6218 856
rect 6386 734 7138 856
rect 7306 734 7966 856
rect 8134 734 8794 856
rect 8962 734 9622 856
rect 9790 734 10542 856
rect 10710 734 11370 856
rect 11538 734 12198 856
rect 12366 734 13026 856
rect 13194 734 13946 856
rect 14114 734 14774 856
rect 14942 734 15602 856
rect 15770 734 16430 856
rect 16598 734 17350 856
rect 17518 734 18178 856
rect 18346 734 19006 856
rect 19174 734 19834 856
rect 20002 734 20754 856
rect 20922 734 21582 856
rect 21750 734 22410 856
rect 22578 734 23330 856
rect 23498 734 24158 856
rect 24326 734 24986 856
rect 25154 734 25814 856
rect 25982 734 26734 856
rect 26902 734 27562 856
rect 27730 734 28390 856
rect 28558 734 29218 856
rect 29386 734 30138 856
rect 30306 734 30966 856
rect 31134 734 31794 856
rect 31962 734 32622 856
rect 32790 734 33542 856
rect 33710 734 34370 856
rect 34538 734 35198 856
rect 35366 734 36026 856
rect 36194 734 36946 856
rect 37114 734 37774 856
rect 37942 734 38602 856
rect 38770 734 39430 856
rect 39598 734 40350 856
rect 40518 734 41178 856
rect 41346 734 42006 856
rect 42174 734 42834 856
rect 43002 734 43754 856
rect 43922 734 44582 856
rect 44750 734 45410 856
rect 45578 734 46330 856
rect 46498 734 47158 856
rect 47326 734 47986 856
rect 48154 734 48814 856
rect 48982 734 49734 856
rect 49902 734 50562 856
rect 50730 734 51390 856
rect 51558 734 52218 856
rect 52386 734 53138 856
rect 53306 734 53966 856
rect 54134 734 54794 856
rect 54962 734 55622 856
rect 55790 734 56542 856
rect 56710 734 57370 856
rect 57538 734 58198 856
rect 58366 734 59026 856
rect 59194 734 59946 856
rect 60114 734 60774 856
rect 60942 734 61602 856
rect 61770 734 62430 856
rect 62598 734 63350 856
rect 63518 734 64178 856
rect 64346 734 65006 856
rect 65174 734 65834 856
rect 66002 734 66754 856
rect 66922 734 67582 856
rect 67750 734 68410 856
rect 68578 734 69330 856
rect 69498 734 70158 856
rect 70326 734 70986 856
rect 71154 734 71814 856
rect 71982 734 72734 856
rect 72902 734 73562 856
rect 73730 734 74390 856
rect 74558 734 75218 856
rect 75386 734 76138 856
rect 76306 734 76966 856
rect 77134 734 77794 856
rect 77962 734 78622 856
rect 78790 734 79542 856
rect 79710 734 80370 856
rect 80538 734 81198 856
rect 81366 734 82026 856
rect 82194 734 82946 856
rect 83114 734 83774 856
rect 83942 734 84602 856
rect 84770 734 85430 856
rect 85598 734 86350 856
rect 86518 734 87178 856
rect 87346 734 88006 856
rect 88174 734 88926 856
rect 89094 734 89754 856
rect 89922 734 90582 856
rect 90750 734 91410 856
rect 91578 734 92330 856
rect 92498 734 93158 856
rect 93326 734 93986 856
rect 94154 734 94814 856
rect 94982 734 95734 856
rect 95902 734 96562 856
rect 96730 734 97390 856
rect 97558 734 98218 856
rect 98386 734 99138 856
rect 99306 734 99966 856
rect 100134 734 100794 856
rect 100962 734 101622 856
rect 101790 734 102542 856
rect 102710 734 103370 856
rect 103538 734 104198 856
rect 104366 734 105026 856
rect 105194 734 105946 856
rect 106114 734 106774 856
rect 106942 734 107602 856
rect 107770 734 108430 856
rect 108598 734 109350 856
rect 109518 734 110178 856
rect 110346 734 111006 856
rect 111174 734 111926 856
rect 112094 734 112754 856
rect 112922 734 113582 856
rect 113750 734 114410 856
rect 114578 734 115330 856
rect 115498 734 116158 856
rect 116326 734 116986 856
rect 117154 734 117814 856
rect 117982 734 118734 856
rect 118902 734 119562 856
rect 119730 734 120390 856
rect 120558 734 121218 856
rect 121386 734 122138 856
rect 122306 734 122966 856
rect 123134 734 123794 856
rect 123962 734 124622 856
rect 124790 734 125542 856
rect 125710 734 126370 856
rect 126538 734 127198 856
rect 127366 734 128026 856
rect 128194 734 128946 856
rect 129114 734 129774 856
rect 129942 734 130602 856
rect 130770 734 131430 856
rect 131598 734 132350 856
rect 132518 734 133178 856
rect 133346 734 134006 856
rect 134174 734 134926 856
rect 135094 734 135754 856
rect 135922 734 136582 856
rect 136750 734 137410 856
rect 137578 734 138330 856
rect 138498 734 139158 856
rect 139326 734 139986 856
rect 140154 734 140814 856
rect 140982 734 141734 856
rect 141902 734 142562 856
rect 142730 734 143390 856
rect 143558 734 144218 856
rect 144386 734 145138 856
rect 145306 734 145966 856
rect 146134 734 146794 856
rect 146962 734 147622 856
rect 147790 734 148542 856
rect 148710 734 149370 856
rect 149538 734 150198 856
rect 150366 734 151026 856
rect 151194 734 151946 856
rect 152114 734 152774 856
rect 152942 734 153602 856
rect 153770 734 154430 856
rect 154598 734 155350 856
rect 155518 734 156178 856
rect 156346 734 157006 856
rect 157174 734 157926 856
rect 158094 734 158754 856
rect 158922 734 159582 856
rect 159750 734 160410 856
rect 160578 734 161330 856
rect 161498 734 162158 856
rect 162326 734 162986 856
rect 163154 734 163814 856
rect 163982 734 164734 856
rect 164902 734 165562 856
rect 165730 734 166390 856
rect 166558 734 167218 856
rect 167386 734 168138 856
rect 168306 734 168966 856
rect 169134 734 169794 856
rect 169962 734 170622 856
rect 170790 734 171542 856
rect 171710 734 172370 856
rect 172538 734 173198 856
rect 173366 734 174026 856
rect 174194 734 174946 856
rect 175114 734 175774 856
rect 175942 734 176602 856
rect 176770 734 177522 856
rect 177690 734 178350 856
rect 178518 734 179178 856
rect 179346 734 180006 856
rect 180174 734 180926 856
rect 181094 734 181754 856
rect 181922 734 182582 856
rect 182750 734 183410 856
rect 183578 734 184330 856
rect 184498 734 185158 856
rect 185326 734 185986 856
rect 186154 734 186814 856
rect 186982 734 187734 856
rect 187902 734 188562 856
rect 188730 734 189390 856
rect 189558 734 190218 856
rect 190386 734 191138 856
rect 191306 734 191966 856
rect 192134 734 192794 856
rect 192962 734 193622 856
rect 193790 734 194542 856
rect 194710 734 195370 856
rect 195538 734 196198 856
rect 196366 734 197026 856
rect 197194 734 197946 856
rect 198114 734 198774 856
rect 198942 734 199602 856
rect 199770 734 200522 856
rect 200690 734 201350 856
rect 201518 734 202178 856
rect 202346 734 203006 856
rect 203174 734 203926 856
rect 204094 734 204754 856
rect 204922 734 205582 856
rect 205750 734 206410 856
rect 206578 734 207330 856
rect 207498 734 208158 856
rect 208326 734 208986 856
rect 209154 734 209814 856
rect 209982 734 210734 856
rect 210902 734 211562 856
rect 211730 734 212390 856
rect 212558 734 213218 856
rect 213386 734 214138 856
rect 214306 734 214966 856
rect 215134 734 215794 856
rect 215962 734 216622 856
rect 216790 734 217542 856
rect 217710 734 218370 856
rect 218538 734 219198 856
rect 219366 734 220026 856
rect 220194 734 220946 856
rect 221114 734 221774 856
rect 221942 734 222602 856
rect 222770 734 223522 856
rect 223690 734 224350 856
rect 224518 734 225178 856
rect 225346 734 226006 856
rect 226174 734 226926 856
rect 227094 734 227754 856
rect 227922 734 228582 856
rect 228750 734 229410 856
rect 229578 734 230330 856
rect 230498 734 231158 856
rect 231326 734 231986 856
rect 232154 734 232814 856
rect 232982 734 233734 856
rect 233902 734 234562 856
rect 234730 734 235390 856
rect 235558 734 236218 856
rect 236386 734 237138 856
rect 237306 734 237966 856
rect 238134 734 238794 856
rect 238962 734 239622 856
rect 239790 734 240542 856
rect 240710 734 241370 856
rect 241538 734 242198 856
rect 242366 734 243026 856
rect 243194 734 243946 856
rect 244114 734 244774 856
rect 244942 734 245602 856
rect 245770 734 246522 856
rect 246690 734 247350 856
rect 247518 734 248178 856
rect 248346 734 249006 856
rect 249174 734 249926 856
rect 250094 734 250754 856
rect 250922 734 251582 856
rect 251750 734 252410 856
rect 252578 734 253330 856
rect 253498 734 254158 856
rect 254326 734 254986 856
rect 255154 734 255814 856
rect 255982 734 256734 856
rect 256902 734 257562 856
rect 257730 734 258390 856
rect 258558 734 259218 856
rect 259386 734 260138 856
rect 260306 734 260966 856
rect 261134 734 261794 856
rect 261962 734 262622 856
rect 262790 734 263542 856
rect 263710 734 264370 856
rect 264538 734 265198 856
rect 265366 734 266118 856
rect 266286 734 266946 856
rect 267114 734 267774 856
rect 267942 734 268602 856
rect 268770 734 269522 856
rect 269690 734 270350 856
rect 270518 734 271178 856
rect 271346 734 272006 856
rect 272174 734 272926 856
rect 273094 734 273754 856
rect 273922 734 274582 856
rect 274750 734 275410 856
rect 275578 734 276330 856
rect 276498 734 277158 856
rect 277326 734 277986 856
rect 278154 734 278814 856
rect 278982 734 279734 856
rect 279902 734 280562 856
rect 280730 734 281390 856
rect 281558 734 282218 856
rect 282386 734 283138 856
rect 283306 734 283966 856
rect 284134 734 284794 856
rect 284962 734 285622 856
rect 285790 734 286542 856
rect 286710 734 287370 856
rect 287538 734 288198 856
rect 288366 734 289118 856
rect 289286 734 289946 856
rect 290114 734 290774 856
rect 290942 734 291602 856
rect 291770 734 292522 856
rect 292690 734 293350 856
rect 293518 734 294178 856
rect 294346 734 295006 856
rect 295174 734 295926 856
rect 296094 734 296754 856
rect 296922 734 297582 856
rect 297750 734 298410 856
rect 298578 734 299330 856
rect 299498 734 300158 856
rect 300326 734 300986 856
rect 301154 734 301814 856
rect 301982 734 302734 856
rect 302902 734 303562 856
rect 303730 734 304390 856
rect 304558 734 305218 856
rect 305386 734 306138 856
rect 306306 734 306966 856
rect 307134 734 307794 856
rect 307962 734 308622 856
rect 308790 734 309542 856
rect 309710 734 310370 856
rect 310538 734 311198 856
rect 311366 734 312118 856
rect 312286 734 312946 856
rect 313114 734 313774 856
rect 313942 734 314602 856
rect 314770 734 315522 856
rect 315690 734 316350 856
rect 316518 734 317178 856
rect 317346 734 318006 856
rect 318174 734 318926 856
rect 319094 734 319754 856
rect 319922 734 320582 856
rect 320750 734 321410 856
rect 321578 734 322330 856
rect 322498 734 323158 856
rect 323326 734 323986 856
rect 324154 734 324814 856
rect 324982 734 325734 856
rect 325902 734 326562 856
rect 326730 734 327390 856
rect 327558 734 328218 856
rect 328386 734 329138 856
rect 329306 734 329966 856
rect 330134 734 330794 856
rect 330962 734 331622 856
rect 331790 734 332542 856
rect 332710 734 333370 856
rect 333538 734 334198 856
rect 334366 734 335118 856
rect 335286 734 335946 856
rect 336114 734 336774 856
rect 336942 734 337602 856
rect 337770 734 338522 856
rect 338690 734 339350 856
rect 339518 734 340178 856
rect 340346 734 341006 856
rect 341174 734 341926 856
rect 342094 734 342754 856
rect 342922 734 343582 856
rect 343750 734 344410 856
rect 344578 734 345330 856
rect 345498 734 346158 856
rect 346326 734 346986 856
rect 347154 734 347814 856
rect 347982 734 348734 856
rect 348902 734 349562 856
rect 349730 734 350390 856
rect 350558 734 351218 856
rect 351386 734 352138 856
rect 352306 734 352966 856
rect 353134 734 353794 856
rect 353962 734 354714 856
rect 354882 734 355542 856
rect 355710 734 356370 856
rect 356538 734 357198 856
rect 357366 734 358118 856
rect 358286 734 358946 856
rect 359114 734 359774 856
rect 359942 734 360602 856
rect 360770 734 361522 856
rect 361690 734 362350 856
rect 362518 734 363178 856
rect 363346 734 364006 856
rect 364174 734 364926 856
rect 365094 734 365754 856
rect 365922 734 366582 856
rect 366750 734 367410 856
rect 367578 734 368330 856
rect 368498 734 369158 856
rect 369326 734 369986 856
rect 370154 734 370814 856
rect 370982 734 371734 856
rect 371902 734 372562 856
rect 372730 734 373390 856
rect 373558 734 374218 856
rect 374386 734 375138 856
rect 375306 734 375966 856
rect 376134 734 376794 856
rect 376962 734 377714 856
rect 377882 734 378542 856
rect 378710 734 379370 856
rect 379538 734 380198 856
rect 380366 734 381118 856
rect 381286 734 381946 856
rect 382114 734 382774 856
rect 382942 734 383602 856
rect 383770 734 384522 856
rect 384690 734 385350 856
rect 385518 734 386178 856
rect 386346 734 387006 856
rect 387174 734 387926 856
rect 388094 734 388754 856
rect 388922 734 389582 856
rect 389750 734 390410 856
rect 390578 734 391330 856
rect 391498 734 392158 856
rect 392326 734 392986 856
rect 393154 734 393814 856
rect 393982 734 394734 856
rect 394902 734 395562 856
rect 395730 734 396390 856
rect 396558 734 397218 856
rect 397386 734 398138 856
rect 398306 734 398966 856
rect 399134 734 399794 856
rect 399962 734 400714 856
rect 400882 734 401542 856
rect 401710 734 402370 856
rect 402538 734 403198 856
rect 403366 734 404118 856
rect 404286 734 404946 856
rect 405114 734 405774 856
rect 405942 734 406602 856
rect 406770 734 407522 856
rect 407690 734 408350 856
rect 408518 734 409178 856
rect 409346 734 410006 856
rect 410174 734 410926 856
rect 411094 734 411754 856
rect 411922 734 412582 856
rect 412750 734 413410 856
rect 413578 734 414330 856
rect 414498 734 415158 856
rect 415326 734 415986 856
rect 416154 734 416814 856
rect 416982 734 417734 856
rect 417902 734 418562 856
rect 418730 734 419390 856
<< obsm3 >>
rect 4208 2143 403888 417825
<< metal4 >>
rect 4208 2128 4528 417840
rect 19568 2128 19888 417840
rect 34928 2128 35248 417840
rect 50288 2128 50608 417840
rect 65648 2128 65968 417840
rect 81008 2128 81328 417840
rect 96368 2128 96688 417840
rect 111728 2128 112048 417840
rect 127088 2128 127408 417840
rect 142448 2128 142768 417840
rect 157808 2128 158128 417840
rect 173168 2128 173488 417840
rect 188528 2128 188848 417840
rect 203888 2128 204208 417840
rect 219248 2128 219568 417840
rect 234608 2128 234928 417840
rect 249968 2128 250288 417840
rect 265328 2128 265648 417840
rect 280688 2128 281008 417840
rect 296048 2128 296368 417840
rect 311408 2128 311728 417840
rect 326768 2128 327088 417840
rect 342128 2128 342448 417840
rect 357488 2128 357808 417840
rect 372848 2128 373168 417840
rect 388208 2128 388528 417840
rect 403568 2128 403888 417840
<< obsm4 >>
rect 87643 23835 96288 274957
rect 96768 23835 111648 274957
rect 112128 23835 127008 274957
rect 127488 23835 142368 274957
rect 142848 23835 157728 274957
rect 158208 23835 173085 274957
<< labels >>
rlabel metal2 s 1858 419200 1914 420000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 112350 419200 112406 420000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 123390 419200 123446 420000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 134430 419200 134486 420000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 145470 419200 145526 420000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 156510 419200 156566 420000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 167550 419200 167606 420000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 178682 419200 178738 420000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 189722 419200 189778 420000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 200762 419200 200818 420000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 211802 419200 211858 420000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 12898 419200 12954 420000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 222842 419200 222898 420000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 233882 419200 233938 420000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 244922 419200 244978 420000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 256054 419200 256110 420000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 267094 419200 267150 420000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 278134 419200 278190 420000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 289174 419200 289230 420000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 300214 419200 300270 420000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 311254 419200 311310 420000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 322294 419200 322350 420000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 23938 419200 23994 420000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 333334 419200 333390 420000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 344466 419200 344522 420000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 355506 419200 355562 420000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 366546 419200 366602 420000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 377586 419200 377642 420000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 388626 419200 388682 420000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 399666 419200 399722 420000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 410706 419200 410762 420000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 34978 419200 35034 420000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 46018 419200 46074 420000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 57058 419200 57114 420000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 68098 419200 68154 420000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 79138 419200 79194 420000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 90270 419200 90326 420000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 101310 419200 101366 420000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5538 419200 5594 420000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 116030 419200 116086 420000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 127070 419200 127126 420000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 138110 419200 138166 420000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 149150 419200 149206 420000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 160190 419200 160246 420000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 171322 419200 171378 420000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 182362 419200 182418 420000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 193402 419200 193458 420000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 204442 419200 204498 420000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 215482 419200 215538 420000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 16578 419200 16634 420000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 226522 419200 226578 420000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 237562 419200 237618 420000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 248602 419200 248658 420000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 259734 419200 259790 420000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 270774 419200 270830 420000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 281814 419200 281870 420000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 292854 419200 292910 420000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 303894 419200 303950 420000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 314934 419200 314990 420000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 325974 419200 326030 420000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 27618 419200 27674 420000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 337014 419200 337070 420000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 348146 419200 348202 420000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 359186 419200 359242 420000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 370226 419200 370282 420000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 381266 419200 381322 420000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 392306 419200 392362 420000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 403346 419200 403402 420000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 414386 419200 414442 420000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 38658 419200 38714 420000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 49698 419200 49754 420000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 60738 419200 60794 420000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 71778 419200 71834 420000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 82818 419200 82874 420000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 93950 419200 94006 420000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 104990 419200 105046 420000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 9218 419200 9274 420000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 119710 419200 119766 420000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 130750 419200 130806 420000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 141790 419200 141846 420000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 152830 419200 152886 420000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 163870 419200 163926 420000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 175002 419200 175058 420000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 186042 419200 186098 420000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 197082 419200 197138 420000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 208122 419200 208178 420000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 219162 419200 219218 420000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 20258 419200 20314 420000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 230202 419200 230258 420000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 241242 419200 241298 420000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 252282 419200 252338 420000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 263414 419200 263470 420000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 274454 419200 274510 420000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 285494 419200 285550 420000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 296534 419200 296590 420000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 307574 419200 307630 420000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 318614 419200 318670 420000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 329654 419200 329710 420000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 31298 419200 31354 420000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 340786 419200 340842 420000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 351826 419200 351882 420000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 362866 419200 362922 420000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 373906 419200 373962 420000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 384946 419200 385002 420000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 395986 419200 396042 420000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 407026 419200 407082 420000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 418066 419200 418122 420000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 42338 419200 42394 420000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 53378 419200 53434 420000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 64418 419200 64474 420000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 75458 419200 75514 420000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 86590 419200 86646 420000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 97630 419200 97686 420000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 108670 419200 108726 420000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 417790 0 417846 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 418618 0 418674 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 419446 0 419502 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 346214 0 346270 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 348790 0 348846 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 351274 0 351330 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 353850 0 353906 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 356426 0 356482 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 359002 0 359058 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 361578 0 361634 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 364062 0 364118 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 366638 0 366694 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 369214 0 369270 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 371790 0 371846 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 374274 0 374330 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 376850 0 376906 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 379426 0 379482 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 382002 0 382058 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 384578 0 384634 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 387062 0 387118 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 389638 0 389694 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 392214 0 392270 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 394790 0 394846 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 397274 0 397330 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 399850 0 399906 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 402426 0 402482 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 405002 0 405058 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 407578 0 407634 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 410062 0 410118 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 412638 0 412694 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 415214 0 415270 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 192850 0 192906 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 200578 0 200634 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 205638 0 205694 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 208214 0 208270 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 210790 0 210846 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 213274 0 213330 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 215850 0 215906 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 218426 0 218482 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 221002 0 221058 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 223578 0 223634 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 228638 0 228694 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 236274 0 236330 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 241426 0 241482 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 246578 0 246634 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 249062 0 249118 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 251638 0 251694 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 254214 0 254270 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 256790 0 256846 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 259274 0 259330 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 261850 0 261906 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 264426 0 264482 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 267002 0 267058 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 269578 0 269634 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 272062 0 272118 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 274638 0 274694 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 277214 0 277270 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 279790 0 279846 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 282274 0 282330 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 284850 0 284906 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 287426 0 287482 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 290002 0 290058 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 292578 0 292634 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 295062 0 295118 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 297638 0 297694 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 300214 0 300270 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 305274 0 305330 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 307850 0 307906 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 310426 0 310482 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 313002 0 313058 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 315578 0 315634 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 318062 0 318118 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 320638 0 320694 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 323214 0 323270 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 325790 0 325846 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 328274 0 328330 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 330850 0 330906 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 333426 0 333482 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 336002 0 336058 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 338578 0 338634 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 341062 0 341118 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 343638 0 343694 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 347042 0 347098 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 349618 0 349674 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 352194 0 352250 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 354770 0 354826 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 357254 0 357310 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 359830 0 359886 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 362406 0 362462 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 364982 0 365038 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 367466 0 367522 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 370042 0 370098 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 372618 0 372674 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 375194 0 375250 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 377770 0 377826 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 380254 0 380310 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 382830 0 382886 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 385406 0 385462 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 387982 0 388038 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 390466 0 390522 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 393042 0 393098 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 395618 0 395674 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 398194 0 398250 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 400770 0 400826 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 403254 0 403310 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 405830 0 405886 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 408406 0 408462 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 410982 0 411038 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 413466 0 413522 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 416042 0 416098 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 140042 0 140098 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 145194 0 145250 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 150254 0 150310 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 152830 0 152886 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 157982 0 158038 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 163042 0 163098 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 168194 0 168250 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 178406 0 178462 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 180982 0 181038 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 183466 0 183522 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 186042 0 186098 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 188618 0 188674 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 191194 0 191250 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 193678 0 193734 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 196254 0 196310 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 198830 0 198886 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 201406 0 201462 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 203982 0 204038 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 206466 0 206522 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 209042 0 209098 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 211618 0 211674 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 214194 0 214250 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 216678 0 216734 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 219254 0 219310 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 221830 0 221886 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 224406 0 224462 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 226982 0 227038 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 229466 0 229522 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 232042 0 232098 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 234618 0 234674 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 237194 0 237250 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 239678 0 239734 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 242254 0 242310 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 244830 0 244886 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 247406 0 247462 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 249982 0 250038 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 252466 0 252522 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 255042 0 255098 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 257618 0 257674 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 260194 0 260250 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 262678 0 262734 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 265254 0 265310 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 267830 0 267886 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 270406 0 270462 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 272982 0 273038 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 275466 0 275522 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 278042 0 278098 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 280618 0 280674 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 283194 0 283250 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 285678 0 285734 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 288254 0 288310 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 290830 0 290886 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 293406 0 293462 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 295982 0 296038 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 298466 0 298522 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 301042 0 301098 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 303618 0 303674 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 306194 0 306250 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 308678 0 308734 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 311254 0 311310 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 313830 0 313886 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 316406 0 316462 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 318982 0 319038 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 321466 0 321522 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 324042 0 324098 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 326618 0 326674 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 329194 0 329250 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 331678 0 331734 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 334254 0 334310 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 336830 0 336886 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 339406 0 339462 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 341982 0 342038 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 344466 0 344522 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 347870 0 347926 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 350446 0 350502 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 353022 0 353078 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 355598 0 355654 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 358174 0 358230 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 360658 0 360714 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 363234 0 363290 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 365810 0 365866 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 368386 0 368442 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 370870 0 370926 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 373446 0 373502 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 376022 0 376078 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 378598 0 378654 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 381174 0 381230 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 383658 0 383714 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 386234 0 386290 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 388810 0 388866 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 391386 0 391442 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 393870 0 393926 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 396446 0 396502 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 399022 0 399078 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 401598 0 401654 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 404174 0 404230 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 406658 0 406714 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 409234 0 409290 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 411810 0 411866 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 414386 0 414442 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 416870 0 416926 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 181810 0 181866 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 184386 0 184442 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 186870 0 186926 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 189446 0 189502 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 194598 0 194654 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 197082 0 197138 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 207386 0 207442 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 212446 0 212502 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 217598 0 217654 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 220082 0 220138 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 225234 0 225290 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 227810 0 227866 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 230386 0 230442 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 232870 0 232926 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 240598 0 240654 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 243082 0 243138 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 245658 0 245714 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 248234 0 248290 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 250810 0 250866 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 255870 0 255926 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 258446 0 258502 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 261022 0 261078 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 266174 0 266230 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 268658 0 268714 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 271234 0 271290 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 273810 0 273866 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 276386 0 276442 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 278870 0 278926 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 281446 0 281502 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 284022 0 284078 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 286598 0 286654 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 289174 0 289230 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 291658 0 291714 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 294234 0 294290 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 296810 0 296866 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 299386 0 299442 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 301870 0 301926 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 304446 0 304502 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 307022 0 307078 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 309598 0 309654 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 312174 0 312230 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 314658 0 314714 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 317234 0 317290 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 319810 0 319866 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 322386 0 322442 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 324870 0 324926 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 327446 0 327502 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 330022 0 330078 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 332598 0 332654 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 335174 0 335230 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 337658 0 337714 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 340234 0 340290 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 342810 0 342866 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 345386 0 345442 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 403568 2128 403888 417840 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 417840 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 417840 6 vssd1
port 503 nsew ground input
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 82082 0 82138 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 420000 420000
string LEFview TRUE
string GDS_FILE /project/openlane/computer/runs/computer/results/magic/computer.gds
string GDS_END 114024662
string GDS_START 956080
<< end >>

