magic
tech sky130A
magscale 1 2
timestamp 1635000722
<< locali >>
rect 170539 701437 170689 701471
rect 170447 701301 170597 701335
rect 170447 701165 170631 701199
rect 170321 700859 170355 701097
rect 170597 701063 170631 701165
rect 202797 700587 202831 701097
rect 257077 700247 257111 701097
rect 267657 700723 267691 701097
rect 283849 700791 283883 701097
rect 300133 700655 300167 701097
rect 304917 700315 304951 701097
rect 330217 700383 330251 701097
rect 332517 700383 332551 701097
rect 342177 700927 342211 701097
rect 345029 700859 345063 701097
rect 345397 700655 345431 700825
rect 345489 700655 345523 701097
rect 348709 700927 348743 701097
rect 351929 700927 351963 701029
rect 351837 700315 351871 700893
rect 352021 700383 352055 701029
rect 354597 700859 354631 701097
rect 356529 700859 356563 701097
rect 359289 701097 359565 701131
rect 359289 701063 359323 701097
rect 367201 700519 367235 702253
rect 367109 700383 367143 700485
rect 352113 700315 352147 700349
rect 351837 700281 352147 700315
rect 367017 700315 367051 700349
rect 367477 700315 367511 701097
rect 378149 700723 378183 701097
rect 381645 700791 381679 701097
rect 389189 700587 389223 701097
rect 396917 701029 397193 701063
rect 396917 700995 396951 701029
rect 397469 700859 397503 701097
rect 403725 700451 403759 701097
rect 367017 700281 367511 700315
rect 411269 700111 411303 701097
rect 414765 700179 414799 701097
rect 422401 699771 422435 701097
rect 425897 699975 425931 701097
rect 433349 699771 433383 701097
rect 436937 700043 436971 701097
rect 444389 699907 444423 701097
rect 455429 699839 455463 701097
rect 462329 700655 462363 701097
rect 254961 279531 254995 279701
rect 317429 279599 317463 279973
rect 324053 279939 324087 280109
rect 255053 279395 255087 279497
rect 324145 279123 324179 280109
rect 325743 279973 326445 280007
rect 519461 279973 519829 280007
rect 519461 279735 519495 279973
rect 335001 279191 335035 279565
rect 359841 279191 359875 279361
rect 410809 278851 410843 279565
rect 425621 279327 425655 279633
rect 469597 278919 469631 279497
rect 527557 279055 527591 279973
rect 582389 10319 582423 701097
rect 582481 126055 582515 702593
rect 582573 45543 582607 701369
rect 582665 59347 582699 701029
rect 582757 71723 582791 701777
rect 582849 85527 582883 701641
rect 582941 245599 582975 702661
rect 40785 3383 40819 4029
rect 228189 3519 228223 4097
rect 239045 3655 239079 4029
rect 38301 3247 38335 3349
rect 85589 3111 85623 3281
rect 118709 2907 118743 3077
rect 164801 2839 164835 3485
rect 238953 3247 238987 3621
rect 239229 3519 239263 4097
rect 286425 3859 286459 4029
rect 325065 3383 325099 3553
rect 298385 3111 298419 3349
rect 326721 3111 326755 3417
rect 354689 3383 354723 3757
rect 298293 2839 298327 3077
rect 302249 2975 302283 3077
rect 355333 2975 355367 3485
rect 383025 2907 383059 3349
rect 392685 2907 392719 3281
rect 396733 3247 396767 4097
rect 421021 3723 421055 3893
rect 424885 3655 424919 3893
rect 437673 3893 437857 3927
rect 437673 3791 437707 3893
rect 447057 3859 447091 3961
rect 447057 3825 447241 3859
rect 399585 2839 399619 3553
rect 404737 2839 404771 3485
rect 415501 3043 415535 3621
rect 419549 3111 419583 3485
rect 423689 3383 423723 3621
rect 415351 3009 415535 3043
rect 433165 2975 433199 3757
rect 437765 3315 437799 3757
rect 443745 3587 443779 3825
rect 435465 2975 435499 3281
rect 440249 2975 440283 3349
rect 450645 3315 450679 3553
rect 451289 3315 451323 3417
rect 465733 3043 465767 4097
rect 501521 3723 501555 3893
rect 471529 3383 471563 3621
rect 489285 3315 489319 3553
rect 501613 3519 501647 3689
rect 583033 3519 583067 279633
<< viali >>
rect 582941 702661 582975 702695
rect 582481 702593 582515 702627
rect 367201 702253 367235 702287
rect 170505 701437 170539 701471
rect 170689 701437 170723 701471
rect 170413 701301 170447 701335
rect 170597 701301 170631 701335
rect 170413 701165 170447 701199
rect 170321 701097 170355 701131
rect 170597 701029 170631 701063
rect 202797 701097 202831 701131
rect 170321 700825 170355 700859
rect 202797 700553 202831 700587
rect 257077 701097 257111 701131
rect 267657 701097 267691 701131
rect 283849 701097 283883 701131
rect 283849 700757 283883 700791
rect 300133 701097 300167 701131
rect 267657 700689 267691 700723
rect 300133 700621 300167 700655
rect 304917 701097 304951 701131
rect 330217 701097 330251 701131
rect 330217 700349 330251 700383
rect 332517 701097 332551 701131
rect 342177 701097 342211 701131
rect 342177 700893 342211 700927
rect 345029 701097 345063 701131
rect 345489 701097 345523 701131
rect 345029 700825 345063 700859
rect 345397 700825 345431 700859
rect 345397 700621 345431 700655
rect 348709 701097 348743 701131
rect 354597 701097 354631 701131
rect 351929 701029 351963 701063
rect 348709 700893 348743 700927
rect 351837 700893 351871 700927
rect 351929 700893 351963 700927
rect 352021 701029 352055 701063
rect 345489 700621 345523 700655
rect 332517 700349 332551 700383
rect 304917 700281 304951 700315
rect 354597 700825 354631 700859
rect 356529 701097 356563 701131
rect 359565 701097 359599 701131
rect 359289 701029 359323 701063
rect 356529 700825 356563 700859
rect 367109 700485 367143 700519
rect 367201 700485 367235 700519
rect 367477 701097 367511 701131
rect 352021 700349 352055 700383
rect 352113 700349 352147 700383
rect 367017 700349 367051 700383
rect 367109 700349 367143 700383
rect 378149 701097 378183 701131
rect 381645 701097 381679 701131
rect 381645 700757 381679 700791
rect 389189 701097 389223 701131
rect 378149 700689 378183 700723
rect 397469 701097 397503 701131
rect 397193 701029 397227 701063
rect 396917 700961 396951 700995
rect 397469 700825 397503 700859
rect 403725 701097 403759 701131
rect 389189 700553 389223 700587
rect 403725 700417 403759 700451
rect 411269 701097 411303 701131
rect 257077 700213 257111 700247
rect 414765 701097 414799 701131
rect 414765 700145 414799 700179
rect 422401 701097 422435 701131
rect 411269 700077 411303 700111
rect 425897 701097 425931 701131
rect 425897 699941 425931 699975
rect 433349 701097 433383 701131
rect 422401 699737 422435 699771
rect 436937 701097 436971 701131
rect 436937 700009 436971 700043
rect 444389 701097 444423 701131
rect 444389 699873 444423 699907
rect 455429 701097 455463 701131
rect 462329 701097 462363 701131
rect 462329 700621 462363 700655
rect 582389 701097 582423 701131
rect 455429 699805 455463 699839
rect 433349 699737 433383 699771
rect 324053 280109 324087 280143
rect 317429 279973 317463 280007
rect 254961 279701 254995 279735
rect 324053 279905 324087 279939
rect 324145 280109 324179 280143
rect 317429 279565 317463 279599
rect 254961 279497 254995 279531
rect 255053 279497 255087 279531
rect 255053 279361 255087 279395
rect 325709 279973 325743 280007
rect 326445 279973 326479 280007
rect 519829 279973 519863 280007
rect 527557 279973 527591 280007
rect 519461 279701 519495 279735
rect 425621 279633 425655 279667
rect 335001 279565 335035 279599
rect 410809 279565 410843 279599
rect 335001 279157 335035 279191
rect 359841 279361 359875 279395
rect 359841 279157 359875 279191
rect 324145 279089 324179 279123
rect 425621 279293 425655 279327
rect 469597 279497 469631 279531
rect 527557 279021 527591 279055
rect 469597 278885 469631 278919
rect 410809 278817 410843 278851
rect 582757 701777 582791 701811
rect 582481 126021 582515 126055
rect 582573 701369 582607 701403
rect 582665 701029 582699 701063
rect 582849 701641 582883 701675
rect 582941 245565 582975 245599
rect 583033 279633 583067 279667
rect 582849 85493 582883 85527
rect 582757 71689 582791 71723
rect 582665 59313 582699 59347
rect 582573 45509 582607 45543
rect 582389 10285 582423 10319
rect 228189 4097 228223 4131
rect 40785 4029 40819 4063
rect 239229 4097 239263 4131
rect 239045 4029 239079 4063
rect 38301 3349 38335 3383
rect 40785 3349 40819 3383
rect 164801 3485 164835 3519
rect 228189 3485 228223 3519
rect 238953 3621 238987 3655
rect 239045 3621 239079 3655
rect 38301 3213 38335 3247
rect 85589 3281 85623 3315
rect 85589 3077 85623 3111
rect 118709 3077 118743 3111
rect 118709 2873 118743 2907
rect 396733 4097 396767 4131
rect 286425 4029 286459 4063
rect 286425 3825 286459 3859
rect 354689 3757 354723 3791
rect 239229 3485 239263 3519
rect 325065 3553 325099 3587
rect 238953 3213 238987 3247
rect 298385 3349 298419 3383
rect 325065 3349 325099 3383
rect 326721 3417 326755 3451
rect 354689 3349 354723 3383
rect 355333 3485 355367 3519
rect 164801 2805 164835 2839
rect 298293 3077 298327 3111
rect 298385 3077 298419 3111
rect 302249 3077 302283 3111
rect 326721 3077 326755 3111
rect 302249 2941 302283 2975
rect 355333 2941 355367 2975
rect 383025 3349 383059 3383
rect 383025 2873 383059 2907
rect 392685 3281 392719 3315
rect 465733 4097 465767 4131
rect 447057 3961 447091 3995
rect 421021 3893 421055 3927
rect 421021 3689 421055 3723
rect 424885 3893 424919 3927
rect 437857 3893 437891 3927
rect 443745 3825 443779 3859
rect 447241 3825 447275 3859
rect 415501 3621 415535 3655
rect 396733 3213 396767 3247
rect 399585 3553 399619 3587
rect 392685 2873 392719 2907
rect 298293 2805 298327 2839
rect 399585 2805 399619 2839
rect 404737 3485 404771 3519
rect 423689 3621 423723 3655
rect 424885 3621 424919 3655
rect 433165 3757 433199 3791
rect 437673 3757 437707 3791
rect 437765 3757 437799 3791
rect 419549 3485 419583 3519
rect 423689 3349 423723 3383
rect 419549 3077 419583 3111
rect 415317 3009 415351 3043
rect 443745 3553 443779 3587
rect 450645 3553 450679 3587
rect 433165 2941 433199 2975
rect 435465 3281 435499 3315
rect 437765 3281 437799 3315
rect 440249 3349 440283 3383
rect 435465 2941 435499 2975
rect 450645 3281 450679 3315
rect 451289 3417 451323 3451
rect 451289 3281 451323 3315
rect 501521 3893 501555 3927
rect 501521 3689 501555 3723
rect 501613 3689 501647 3723
rect 471529 3621 471563 3655
rect 471529 3349 471563 3383
rect 489285 3553 489319 3587
rect 501613 3485 501647 3519
rect 583033 3485 583067 3519
rect 489285 3281 489319 3315
rect 465733 3009 465767 3043
rect 440249 2941 440283 2975
rect 404737 2805 404771 2839
<< metal1 >>
rect 141418 703604 141424 703656
rect 141476 703644 141482 703656
rect 551094 703644 551100 703656
rect 141476 703616 551100 703644
rect 141476 703604 141482 703616
rect 551094 703604 551100 703616
rect 551152 703604 551158 703656
rect 345014 703536 345020 703588
rect 345072 703576 345078 703588
rect 396350 703576 396356 703588
rect 345072 703548 396356 703576
rect 345072 703536 345078 703548
rect 396350 703536 396356 703548
rect 396408 703536 396414 703588
rect 342162 703468 342168 703520
rect 342220 703508 342226 703520
rect 407390 703508 407396 703520
rect 342220 703480 407396 703508
rect 342220 703468 342226 703480
rect 407390 703468 407396 703480
rect 407448 703468 407454 703520
rect 275462 703400 275468 703452
rect 275520 703440 275526 703452
rect 351178 703440 351184 703452
rect 275520 703412 351184 703440
rect 275520 703400 275526 703412
rect 351178 703400 351184 703412
rect 351236 703400 351242 703452
rect 352834 703400 352840 703452
rect 352892 703440 352898 703452
rect 429838 703440 429844 703452
rect 352892 703412 429844 703440
rect 352892 703400 352898 703412
rect 429838 703400 429844 703412
rect 429896 703400 429902 703452
rect 161566 703332 161572 703384
rect 161624 703372 161630 703384
rect 346394 703372 346400 703384
rect 161624 703344 346400 703372
rect 161624 703332 161630 703344
rect 346394 703332 346400 703344
rect 346452 703332 346458 703384
rect 349062 703332 349068 703384
rect 349120 703372 349126 703384
rect 478506 703372 478512 703384
rect 349120 703344 478512 703372
rect 349120 703332 349126 703344
rect 478506 703332 478512 703344
rect 478564 703332 478570 703384
rect 235166 703264 235172 703316
rect 235224 703304 235230 703316
rect 385310 703304 385316 703316
rect 235224 703276 385316 703304
rect 235224 703264 235230 703276
rect 385310 703264 385316 703276
rect 385368 703264 385374 703316
rect 340414 703196 340420 703248
rect 340472 703236 340478 703248
rect 577038 703236 577044 703248
rect 340472 703208 577044 703236
rect 340472 703196 340478 703208
rect 577038 703196 577044 703208
rect 577096 703196 577102 703248
rect 164786 703128 164792 703180
rect 164844 703168 164850 703180
rect 440602 703168 440608 703180
rect 164844 703140 440608 703168
rect 164844 703128 164850 703140
rect 440602 703128 440608 703140
rect 440660 703128 440666 703180
rect 164510 703060 164516 703112
rect 164568 703100 164574 703112
rect 451642 703100 451648 703112
rect 164568 703072 451648 703100
rect 164568 703060 164574 703072
rect 451642 703060 451648 703072
rect 451700 703060 451706 703112
rect 282822 702992 282828 703044
rect 282880 703032 282886 703044
rect 576946 703032 576952 703044
rect 282880 703004 576952 703032
rect 282880 702992 282886 703004
rect 576946 702992 576952 703004
rect 577004 702992 577010 703044
rect 165338 702924 165344 702976
rect 165396 702964 165402 702976
rect 462682 702964 462688 702976
rect 165396 702936 462688 702964
rect 165396 702924 165402 702936
rect 462682 702924 462688 702936
rect 462740 702924 462746 702976
rect 165154 702856 165160 702908
rect 165212 702896 165218 702908
rect 473722 702896 473728 702908
rect 165212 702868 473728 702896
rect 165212 702856 165218 702868
rect 473722 702856 473728 702868
rect 473780 702856 473786 702908
rect 161842 702788 161848 702840
rect 161900 702828 161906 702840
rect 484762 702828 484768 702840
rect 161900 702800 484768 702828
rect 161900 702788 161906 702800
rect 484762 702788 484768 702800
rect 484820 702788 484826 702840
rect 162026 702720 162032 702772
rect 162084 702760 162090 702772
rect 495802 702760 495808 702772
rect 162084 702732 495808 702760
rect 162084 702720 162090 702732
rect 495802 702720 495808 702732
rect 495860 702720 495866 702772
rect 231210 702652 231216 702704
rect 231268 702692 231274 702704
rect 582929 702695 582987 702701
rect 582929 702692 582941 702695
rect 231268 702664 582941 702692
rect 231268 702652 231274 702664
rect 582929 702661 582941 702664
rect 582975 702661 582987 702695
rect 582929 702655 582987 702661
rect 198090 702584 198096 702636
rect 198148 702624 198154 702636
rect 582469 702627 582527 702633
rect 582469 702624 582481 702627
rect 198148 702596 582481 702624
rect 198148 702584 198154 702596
rect 582469 702593 582481 702596
rect 582515 702593 582527 702627
rect 582469 702587 582527 702593
rect 148318 702516 148324 702568
rect 148376 702556 148382 702568
rect 540054 702556 540060 702568
rect 148376 702528 540060 702556
rect 148376 702516 148382 702528
rect 540054 702516 540060 702528
rect 540112 702516 540118 702568
rect 356054 702448 356060 702500
rect 356112 702488 356118 702500
rect 374270 702488 374276 702500
rect 356112 702460 374276 702488
rect 356112 702448 356118 702460
rect 374270 702448 374276 702460
rect 374328 702448 374334 702500
rect 14458 702380 14464 702432
rect 14516 702420 14522 702432
rect 466454 702420 466460 702432
rect 14516 702392 466460 702420
rect 14516 702380 14522 702392
rect 466454 702380 466460 702392
rect 466512 702380 466518 702432
rect 17218 702312 17224 702364
rect 17276 702352 17282 702364
rect 477494 702352 477500 702364
rect 17276 702324 477500 702352
rect 17276 702312 17282 702324
rect 477494 702312 477500 702324
rect 477552 702312 477558 702364
rect 341794 702244 341800 702296
rect 341852 702284 341858 702296
rect 350442 702284 350448 702296
rect 341852 702256 350448 702284
rect 341852 702244 341858 702256
rect 350442 702244 350448 702256
rect 350500 702244 350506 702296
rect 351178 702244 351184 702296
rect 351236 702284 351242 702296
rect 362494 702284 362500 702296
rect 351236 702256 362500 702284
rect 351236 702244 351242 702256
rect 362494 702244 362500 702256
rect 362552 702244 362558 702296
rect 363874 702244 363880 702296
rect 363932 702284 363938 702296
rect 364978 702284 364984 702296
rect 363932 702256 364984 702284
rect 363932 702244 363938 702256
rect 364978 702244 364984 702256
rect 365036 702244 365042 702296
rect 367186 702284 367192 702296
rect 367147 702256 367192 702284
rect 367186 702244 367192 702256
rect 367244 702244 367250 702296
rect 323302 702176 323308 702228
rect 323360 702216 323366 702228
rect 419350 702216 419356 702228
rect 323360 702188 419356 702216
rect 323360 702176 323366 702188
rect 419350 702176 419356 702188
rect 419408 702176 419414 702228
rect 253382 702108 253388 702160
rect 253440 702148 253446 702160
rect 340414 702148 340420 702160
rect 253440 702120 340420 702148
rect 253440 702108 253446 702120
rect 340414 702108 340420 702120
rect 340472 702108 340478 702160
rect 346394 702108 346400 702160
rect 346452 702148 346458 702160
rect 447962 702148 447968 702160
rect 346452 702120 447968 702148
rect 346452 702108 346458 702120
rect 447962 702108 447968 702120
rect 448020 702108 448026 702160
rect 71038 702040 71044 702092
rect 71096 702080 71102 702092
rect 358722 702080 358728 702092
rect 71096 702052 358728 702080
rect 71096 702040 71102 702052
rect 358722 702040 358728 702052
rect 358780 702040 358786 702092
rect 360286 702080 360292 702092
rect 359016 702052 360292 702080
rect 65518 701972 65524 702024
rect 65576 702012 65582 702024
rect 359016 702012 359044 702052
rect 360286 702040 360292 702052
rect 360344 702040 360350 702092
rect 392670 702080 392676 702092
rect 361684 702052 392676 702080
rect 65576 701984 359044 702012
rect 65576 701972 65582 701984
rect 359090 701972 359096 702024
rect 359148 702012 359154 702024
rect 361684 702012 361712 702052
rect 392670 702040 392676 702052
rect 392728 702040 392734 702092
rect 359148 701984 361712 702012
rect 359148 701972 359154 701984
rect 361758 701972 361764 702024
rect 361816 702012 361822 702024
rect 547414 702012 547420 702024
rect 361816 701984 547420 702012
rect 361816 701972 361822 701984
rect 547414 701972 547420 701984
rect 547472 701972 547478 702024
rect 293540 701904 293546 701956
rect 293598 701944 293604 701956
rect 583478 701944 583484 701956
rect 293598 701916 583484 701944
rect 293598 701904 293604 701916
rect 583478 701904 583484 701916
rect 583536 701904 583542 701956
rect 289860 701836 289866 701888
rect 289918 701876 289924 701888
rect 583570 701876 583576 701888
rect 289918 701848 583576 701876
rect 289918 701836 289924 701848
rect 583570 701836 583576 701848
rect 583628 701836 583634 701888
rect 161658 701768 161664 701820
rect 161716 701808 161722 701820
rect 459002 701808 459008 701820
rect 161716 701780 459008 701808
rect 161716 701768 161722 701780
rect 459002 701768 459008 701780
rect 459060 701768 459066 701820
rect 562778 701768 562784 701820
rect 562836 701808 562842 701820
rect 582745 701811 582803 701817
rect 582745 701808 582757 701811
rect 562836 701780 582757 701808
rect 562836 701768 562842 701780
rect 582745 701777 582757 701780
rect 582791 701777 582803 701811
rect 582745 701771 582803 701777
rect 279142 701700 279148 701752
rect 279200 701740 279206 701752
rect 583386 701740 583392 701752
rect 279200 701712 583392 701740
rect 279200 701700 279206 701712
rect 583386 701700 583392 701712
rect 583444 701700 583450 701752
rect 161750 701632 161756 701684
rect 161808 701672 161814 701684
rect 470042 701672 470048 701684
rect 161808 701644 470048 701672
rect 161808 701632 161814 701644
rect 470042 701632 470048 701644
rect 470100 701632 470106 701684
rect 555418 701632 555424 701684
rect 555476 701672 555482 701684
rect 582837 701675 582895 701681
rect 582837 701672 582849 701675
rect 555476 701644 582849 701672
rect 555476 701632 555482 701644
rect 582837 701641 582849 701644
rect 582883 701641 582895 701675
rect 582837 701635 582895 701641
rect 162118 701564 162124 701616
rect 162176 701604 162182 701616
rect 162176 701576 171134 701604
rect 162176 701564 162182 701576
rect 161934 701496 161940 701548
rect 161992 701536 161998 701548
rect 171106 701536 171134 701576
rect 271782 701564 271788 701616
rect 271840 701604 271846 701616
rect 583202 701604 583208 701616
rect 271840 701576 583208 701604
rect 271840 701564 271846 701576
rect 583202 701564 583208 701576
rect 583260 701564 583266 701616
rect 179046 701536 179052 701548
rect 161992 701508 170628 701536
rect 171106 701508 179052 701536
rect 161992 701496 161998 701508
rect 162394 701428 162400 701480
rect 162452 701468 162458 701480
rect 170493 701471 170551 701477
rect 170493 701468 170505 701471
rect 162452 701440 170505 701468
rect 162452 701428 162458 701440
rect 170493 701437 170505 701440
rect 170539 701437 170551 701471
rect 170493 701431 170551 701437
rect 162210 701360 162216 701412
rect 162268 701400 162274 701412
rect 170600 701400 170628 701508
rect 179046 701496 179052 701508
rect 179104 701496 179110 701548
rect 268102 701496 268108 701548
rect 268160 701536 268166 701548
rect 583294 701536 583300 701548
rect 268160 701508 583300 701536
rect 268160 701496 268166 701508
rect 583294 701496 583300 701508
rect 583352 701496 583358 701548
rect 170677 701471 170735 701477
rect 170677 701437 170689 701471
rect 170723 701468 170735 701471
rect 190086 701468 190092 701480
rect 170723 701440 190092 701468
rect 170723 701437 170735 701440
rect 170677 701431 170735 701437
rect 190086 701428 190092 701440
rect 190144 701428 190150 701480
rect 260742 701428 260748 701480
rect 260800 701468 260806 701480
rect 583018 701468 583024 701480
rect 260800 701440 583024 701468
rect 260800 701428 260806 701440
rect 583018 701428 583024 701440
rect 583076 701428 583082 701480
rect 492122 701400 492128 701412
rect 162268 701372 170536 701400
rect 170600 701372 492128 701400
rect 162268 701360 162274 701372
rect 162486 701292 162492 701344
rect 162544 701332 162550 701344
rect 170401 701335 170459 701341
rect 170401 701332 170413 701335
rect 162544 701304 170413 701332
rect 162544 701292 162550 701304
rect 170401 701301 170413 701304
rect 170447 701301 170459 701335
rect 170401 701295 170459 701301
rect 162302 701224 162308 701276
rect 162360 701264 162366 701276
rect 170508 701264 170536 701372
rect 492122 701360 492128 701372
rect 492180 701360 492186 701412
rect 566458 701360 566464 701412
rect 566516 701400 566522 701412
rect 582561 701403 582619 701409
rect 582561 701400 582573 701403
rect 566516 701372 582573 701400
rect 566516 701360 566522 701372
rect 582561 701369 582573 701372
rect 582607 701369 582619 701403
rect 582561 701363 582619 701369
rect 170585 701335 170643 701341
rect 170585 701301 170597 701335
rect 170631 701332 170643 701335
rect 182726 701332 182732 701344
rect 170631 701304 182732 701332
rect 170631 701301 170643 701304
rect 170585 701295 170643 701301
rect 182726 701292 182732 701304
rect 182784 701292 182790 701344
rect 249702 701292 249708 701344
rect 249760 701332 249766 701344
rect 582834 701332 582840 701344
rect 249760 701304 582840 701332
rect 249760 701292 249766 701304
rect 582834 701292 582840 701304
rect 582892 701292 582898 701344
rect 186406 701264 186412 701276
rect 162360 701236 170444 701264
rect 170508 701236 186412 701264
rect 162360 701224 162366 701236
rect 162578 701156 162584 701208
rect 162636 701196 162642 701208
rect 168006 701196 168012 701208
rect 162636 701168 168012 701196
rect 162636 701156 162642 701168
rect 168006 701156 168012 701168
rect 168064 701156 168070 701208
rect 170416 701205 170444 701236
rect 186406 701224 186412 701236
rect 186464 701224 186470 701276
rect 245746 701224 245752 701276
rect 245804 701264 245810 701276
rect 582926 701264 582932 701276
rect 245804 701236 582932 701264
rect 245804 701224 245810 701236
rect 582926 701224 582932 701236
rect 582984 701224 582990 701276
rect 170401 701199 170459 701205
rect 170401 701165 170413 701199
rect 170447 701165 170459 701199
rect 171686 701196 171692 701208
rect 170401 701159 170459 701165
rect 170508 701168 171692 701196
rect 162762 701088 162768 701140
rect 162820 701128 162826 701140
rect 164326 701128 164332 701140
rect 162820 701100 164332 701128
rect 162820 701088 162826 701100
rect 164326 701088 164332 701100
rect 164384 701088 164390 701140
rect 170306 701128 170312 701140
rect 170267 701100 170312 701128
rect 170306 701088 170312 701100
rect 170364 701088 170370 701140
rect 162670 701020 162676 701072
rect 162728 701060 162734 701072
rect 170508 701060 170536 701168
rect 171686 701156 171692 701168
rect 171744 701156 171750 701208
rect 242250 701156 242256 701208
rect 242308 701196 242314 701208
rect 583754 701196 583760 701208
rect 242308 701168 583760 701196
rect 242308 701156 242314 701168
rect 583754 701156 583760 701168
rect 583812 701156 583818 701208
rect 175366 701128 175372 701140
rect 171106 701100 175372 701128
rect 162728 701032 170536 701060
rect 170585 701063 170643 701069
rect 162728 701020 162734 701032
rect 170585 701029 170597 701063
rect 170631 701060 170643 701063
rect 171106 701060 171134 701100
rect 175366 701088 175372 701100
rect 175424 701088 175430 701140
rect 202782 701128 202788 701140
rect 202743 701100 202788 701128
rect 202782 701088 202788 701100
rect 202840 701088 202846 701140
rect 257062 701128 257068 701140
rect 257023 701100 257068 701128
rect 257062 701088 257068 701100
rect 257120 701088 257126 701140
rect 267642 701128 267648 701140
rect 267603 701100 267648 701128
rect 267642 701088 267648 701100
rect 267700 701088 267706 701140
rect 283834 701128 283840 701140
rect 283795 701100 283840 701128
rect 283834 701088 283840 701100
rect 283892 701088 283898 701140
rect 300118 701128 300124 701140
rect 300079 701100 300124 701128
rect 300118 701088 300124 701100
rect 300176 701088 300182 701140
rect 304902 701128 304908 701140
rect 304863 701100 304908 701128
rect 304902 701088 304908 701100
rect 304960 701088 304966 701140
rect 330202 701128 330208 701140
rect 330163 701100 330208 701128
rect 330202 701088 330208 701100
rect 330260 701088 330266 701140
rect 332502 701128 332508 701140
rect 332463 701100 332508 701128
rect 332502 701088 332508 701100
rect 332560 701088 332566 701140
rect 338022 701088 338028 701140
rect 338080 701088 338086 701140
rect 342162 701128 342168 701140
rect 342123 701100 342168 701128
rect 342162 701088 342168 701100
rect 342220 701088 342226 701140
rect 345014 701088 345020 701140
rect 345072 701128 345078 701140
rect 345474 701128 345480 701140
rect 345072 701100 345117 701128
rect 345435 701100 345480 701128
rect 345072 701088 345078 701100
rect 345474 701088 345480 701100
rect 345532 701088 345538 701140
rect 348694 701128 348700 701140
rect 348655 701100 348700 701128
rect 348694 701088 348700 701100
rect 348752 701088 348758 701140
rect 354585 701131 354643 701137
rect 354585 701097 354597 701131
rect 354631 701128 354643 701131
rect 356054 701128 356060 701140
rect 354631 701100 356060 701128
rect 354631 701097 354643 701100
rect 354585 701091 354643 701097
rect 356054 701088 356060 701100
rect 356112 701088 356118 701140
rect 356514 701128 356520 701140
rect 356475 701100 356520 701128
rect 356514 701088 356520 701100
rect 356572 701088 356578 701140
rect 359458 701088 359464 701140
rect 359516 701088 359522 701140
rect 359553 701131 359611 701137
rect 359553 701097 359565 701131
rect 359599 701128 359611 701131
rect 367094 701128 367100 701140
rect 359599 701100 367100 701128
rect 359599 701097 359611 701100
rect 359553 701091 359611 701097
rect 367094 701088 367100 701100
rect 367152 701088 367158 701140
rect 367465 701131 367523 701137
rect 367465 701097 367477 701131
rect 367511 701128 367523 701131
rect 370590 701128 370596 701140
rect 367511 701100 370596 701128
rect 367511 701097 367523 701100
rect 367465 701091 367523 701097
rect 370590 701088 370596 701100
rect 370648 701088 370654 701140
rect 378134 701128 378140 701140
rect 378095 701100 378140 701128
rect 378134 701088 378140 701100
rect 378192 701088 378198 701140
rect 381630 701128 381636 701140
rect 381591 701100 381636 701128
rect 381630 701088 381636 701100
rect 381688 701088 381694 701140
rect 389174 701128 389180 701140
rect 389135 701100 389180 701128
rect 389174 701088 389180 701100
rect 389232 701088 389238 701140
rect 397454 701128 397460 701140
rect 397415 701100 397460 701128
rect 397454 701088 397460 701100
rect 397512 701088 397518 701140
rect 400214 701088 400220 701140
rect 400272 701088 400278 701140
rect 403710 701128 403716 701140
rect 403671 701100 403716 701128
rect 403710 701088 403716 701100
rect 403768 701088 403774 701140
rect 411254 701128 411260 701140
rect 411215 701100 411260 701128
rect 411254 701088 411260 701100
rect 411312 701088 411318 701140
rect 413646 701088 413652 701140
rect 413704 701088 413710 701140
rect 414750 701128 414756 701140
rect 414711 701100 414756 701128
rect 414750 701088 414756 701100
rect 414808 701088 414814 701140
rect 422386 701128 422392 701140
rect 422347 701100 422392 701128
rect 422386 701088 422392 701100
rect 422444 701088 422450 701140
rect 425882 701128 425888 701140
rect 425843 701100 425888 701128
rect 425882 701088 425888 701100
rect 425940 701088 425946 701140
rect 433334 701128 433340 701140
rect 433295 701100 433340 701128
rect 433334 701088 433340 701100
rect 433392 701088 433398 701140
rect 436922 701128 436928 701140
rect 436883 701100 436928 701128
rect 436922 701088 436928 701100
rect 436980 701088 436986 701140
rect 444374 701128 444380 701140
rect 444335 701100 444380 701128
rect 444374 701088 444380 701100
rect 444432 701088 444438 701140
rect 455414 701128 455420 701140
rect 455375 701100 455420 701128
rect 455414 701088 455420 701100
rect 455472 701088 455478 701140
rect 462314 701128 462320 701140
rect 462275 701100 462320 701128
rect 462314 701088 462320 701100
rect 462372 701088 462378 701140
rect 543458 701088 543464 701140
rect 543516 701088 543522 701140
rect 543734 701088 543740 701140
rect 543792 701088 543798 701140
rect 558454 701088 558460 701140
rect 558512 701088 558518 701140
rect 569954 701088 569960 701140
rect 570012 701128 570018 701140
rect 570012 701100 576854 701128
rect 570012 701088 570018 701100
rect 170631 701032 171134 701060
rect 338040 701060 338068 701088
rect 351917 701063 351975 701069
rect 351917 701060 351929 701063
rect 338040 701032 351929 701060
rect 170631 701029 170643 701032
rect 170585 701023 170643 701029
rect 351917 701029 351929 701032
rect 351963 701029 351975 701063
rect 351917 701023 351975 701029
rect 352009 701063 352067 701069
rect 352009 701029 352021 701063
rect 352055 701060 352067 701063
rect 359277 701063 359335 701069
rect 359277 701060 359289 701063
rect 352055 701032 359289 701060
rect 352055 701029 352067 701032
rect 352009 701023 352067 701029
rect 359277 701029 359289 701032
rect 359323 701029 359335 701063
rect 359476 701060 359504 701088
rect 397181 701063 397239 701069
rect 359476 701032 397132 701060
rect 359277 701023 359335 701029
rect 137830 700952 137836 701004
rect 137888 700992 137894 701004
rect 396905 700995 396963 701001
rect 396905 700992 396917 700995
rect 137888 700964 396917 700992
rect 137888 700952 137894 700964
rect 396905 700961 396917 700964
rect 396951 700961 396963 700995
rect 397104 700992 397132 701032
rect 397181 701029 397193 701063
rect 397227 701060 397239 701063
rect 400232 701060 400260 701088
rect 397227 701032 400260 701060
rect 397227 701029 397239 701032
rect 397181 701023 397239 701029
rect 413664 700992 413692 701088
rect 397104 700964 413692 700992
rect 396905 700955 396963 700961
rect 105446 700884 105452 700936
rect 105504 700924 105510 700936
rect 342165 700927 342223 700933
rect 342165 700924 342177 700927
rect 105504 700896 342177 700924
rect 105504 700884 105510 700896
rect 342165 700893 342177 700896
rect 342211 700893 342223 700927
rect 342165 700887 342223 700893
rect 348697 700927 348755 700933
rect 348697 700893 348709 700927
rect 348743 700924 348755 700927
rect 351825 700927 351883 700933
rect 351825 700924 351837 700927
rect 348743 700896 351837 700924
rect 348743 700893 348755 700896
rect 348697 700887 348755 700893
rect 351825 700893 351837 700896
rect 351871 700893 351883 700927
rect 351825 700887 351883 700893
rect 351917 700927 351975 700933
rect 351917 700893 351929 700927
rect 351963 700924 351975 700927
rect 543476 700924 543504 701088
rect 351963 700896 543504 700924
rect 351963 700893 351975 700896
rect 351917 700887 351975 700893
rect 170309 700859 170367 700865
rect 170309 700825 170321 700859
rect 170355 700856 170367 700859
rect 345017 700859 345075 700865
rect 345017 700856 345029 700859
rect 170355 700828 345029 700856
rect 170355 700825 170367 700828
rect 170309 700819 170367 700825
rect 345017 700825 345029 700828
rect 345063 700825 345075 700859
rect 345017 700819 345075 700825
rect 345385 700859 345443 700865
rect 345385 700825 345397 700859
rect 345431 700856 345443 700859
rect 354585 700859 354643 700865
rect 354585 700856 354597 700859
rect 345431 700828 354597 700856
rect 345431 700825 345443 700828
rect 345385 700819 345443 700825
rect 354585 700825 354597 700828
rect 354631 700825 354643 700859
rect 354585 700819 354643 700825
rect 356517 700859 356575 700865
rect 356517 700825 356529 700859
rect 356563 700856 356575 700859
rect 397457 700859 397515 700865
rect 397457 700856 397469 700859
rect 356563 700828 397469 700856
rect 356563 700825 356575 700828
rect 356517 700819 356575 700825
rect 397457 700825 397469 700828
rect 397503 700825 397515 700859
rect 397457 700819 397515 700825
rect 283837 700791 283895 700797
rect 283837 700757 283849 700791
rect 283883 700788 283895 700791
rect 381633 700791 381691 700797
rect 381633 700788 381645 700791
rect 283883 700760 381645 700788
rect 283883 700757 283895 700760
rect 283837 700751 283895 700757
rect 381633 700757 381645 700760
rect 381679 700757 381691 700791
rect 381633 700751 381691 700757
rect 267645 700723 267703 700729
rect 267645 700689 267657 700723
rect 267691 700720 267703 700723
rect 378137 700723 378195 700729
rect 378137 700720 378149 700723
rect 267691 700692 378149 700720
rect 267691 700689 267703 700692
rect 267645 700683 267703 700689
rect 378137 700689 378149 700692
rect 378183 700689 378195 700723
rect 378137 700683 378195 700689
rect 300121 700655 300179 700661
rect 300121 700621 300133 700655
rect 300167 700652 300179 700655
rect 345385 700655 345443 700661
rect 345385 700652 345397 700655
rect 300167 700624 345397 700652
rect 300167 700621 300179 700624
rect 300121 700615 300179 700621
rect 345385 700621 345397 700624
rect 345431 700621 345443 700655
rect 345385 700615 345443 700621
rect 345477 700655 345535 700661
rect 345477 700621 345489 700655
rect 345523 700652 345535 700655
rect 462317 700655 462375 700661
rect 462317 700652 462329 700655
rect 345523 700624 462329 700652
rect 345523 700621 345535 700624
rect 345477 700615 345535 700621
rect 462317 700621 462329 700624
rect 462363 700621 462375 700655
rect 462317 700615 462375 700621
rect 202785 700587 202843 700593
rect 202785 700553 202797 700587
rect 202831 700584 202843 700587
rect 389177 700587 389235 700593
rect 389177 700584 389189 700587
rect 202831 700556 389189 700584
rect 202831 700553 202843 700556
rect 202785 700547 202843 700553
rect 389177 700553 389189 700556
rect 389223 700553 389235 700587
rect 389177 700547 389235 700553
rect 53098 700476 53104 700528
rect 53156 700516 53162 700528
rect 367097 700519 367155 700525
rect 367097 700516 367109 700519
rect 53156 700488 367109 700516
rect 53156 700476 53162 700488
rect 367097 700485 367109 700488
rect 367143 700485 367155 700519
rect 367097 700479 367155 700485
rect 367189 700519 367247 700525
rect 367189 700485 367201 700519
rect 367235 700516 367247 700519
rect 543752 700516 543780 701088
rect 367235 700488 543780 700516
rect 367235 700485 367247 700488
rect 367189 700479 367247 700485
rect 154114 700408 154120 700460
rect 154172 700448 154178 700460
rect 403713 700451 403771 700457
rect 403713 700448 403725 700451
rect 154172 700420 403725 700448
rect 154172 700408 154178 700420
rect 403713 700417 403725 700420
rect 403759 700417 403771 700451
rect 403713 700411 403771 700417
rect 3418 700340 3424 700392
rect 3476 700380 3482 700392
rect 330205 700383 330263 700389
rect 330205 700380 330217 700383
rect 3476 700352 330217 700380
rect 3476 700340 3482 700352
rect 330205 700349 330217 700352
rect 330251 700349 330263 700383
rect 330205 700343 330263 700349
rect 332505 700383 332563 700389
rect 332505 700349 332517 700383
rect 332551 700380 332563 700383
rect 352009 700383 352067 700389
rect 352009 700380 352021 700383
rect 332551 700352 352021 700380
rect 332551 700349 332563 700352
rect 332505 700343 332563 700349
rect 352009 700349 352021 700352
rect 352055 700349 352067 700383
rect 352009 700343 352067 700349
rect 352101 700383 352159 700389
rect 352101 700349 352113 700383
rect 352147 700380 352159 700383
rect 367005 700383 367063 700389
rect 367005 700380 367017 700383
rect 352147 700352 367017 700380
rect 352147 700349 352159 700352
rect 352101 700343 352159 700349
rect 367005 700349 367017 700352
rect 367051 700349 367063 700383
rect 367005 700343 367063 700349
rect 367097 700383 367155 700389
rect 367097 700349 367109 700383
rect 367143 700380 367155 700383
rect 558472 700380 558500 701088
rect 576826 701060 576854 701100
rect 577498 701088 577504 701140
rect 577556 701128 577562 701140
rect 582377 701131 582435 701137
rect 582377 701128 582389 701131
rect 577556 701100 582389 701128
rect 577556 701088 577562 701100
rect 582377 701097 582389 701100
rect 582423 701097 582435 701131
rect 582377 701091 582435 701097
rect 582653 701063 582711 701069
rect 582653 701060 582665 701063
rect 576826 701032 582665 701060
rect 582653 701029 582665 701032
rect 582699 701029 582711 701063
rect 582653 701023 582711 701029
rect 367143 700352 558500 700380
rect 367143 700349 367155 700352
rect 367097 700343 367155 700349
rect 304905 700315 304963 700321
rect 304905 700281 304917 700315
rect 304951 700312 304963 700315
rect 583662 700312 583668 700324
rect 304951 700284 583668 700312
rect 304951 700281 304963 700284
rect 304905 700275 304963 700281
rect 583662 700272 583668 700284
rect 583720 700272 583726 700324
rect 257065 700247 257123 700253
rect 257065 700213 257077 700247
rect 257111 700244 257123 700247
rect 583110 700244 583116 700256
rect 257111 700216 583116 700244
rect 257111 700213 257123 700216
rect 257065 700207 257123 700213
rect 583110 700204 583116 700216
rect 583168 700204 583174 700256
rect 89162 700136 89168 700188
rect 89220 700176 89226 700188
rect 414753 700179 414811 700185
rect 414753 700176 414765 700179
rect 89220 700148 414765 700176
rect 89220 700136 89226 700148
rect 414753 700145 414765 700148
rect 414799 700145 414811 700179
rect 414753 700139 414811 700145
rect 72970 700068 72976 700120
rect 73028 700108 73034 700120
rect 411257 700111 411315 700117
rect 411257 700108 411269 700111
rect 73028 700080 411269 700108
rect 73028 700068 73034 700080
rect 411257 700077 411269 700080
rect 411303 700077 411315 700111
rect 411257 700071 411315 700077
rect 35158 700000 35164 700052
rect 35216 700040 35222 700052
rect 436925 700043 436983 700049
rect 436925 700040 436937 700043
rect 35216 700012 436937 700040
rect 35216 700000 35222 700012
rect 436925 700009 436937 700012
rect 436971 700009 436983 700043
rect 436925 700003 436983 700009
rect 24302 699932 24308 699984
rect 24360 699972 24366 699984
rect 425885 699975 425943 699981
rect 425885 699972 425897 699975
rect 24360 699944 425897 699972
rect 24360 699932 24366 699944
rect 425885 699941 425897 699944
rect 425931 699941 425943 699975
rect 425885 699935 425943 699941
rect 40678 699864 40684 699916
rect 40736 699904 40742 699916
rect 444377 699907 444435 699913
rect 444377 699904 444389 699907
rect 40736 699876 444389 699904
rect 40736 699864 40742 699876
rect 444377 699873 444389 699876
rect 444423 699873 444435 699907
rect 444377 699867 444435 699873
rect 43438 699796 43444 699848
rect 43496 699836 43502 699848
rect 455417 699839 455475 699845
rect 455417 699836 455429 699839
rect 43496 699808 455429 699836
rect 43496 699796 43502 699808
rect 455417 699805 455429 699808
rect 455463 699805 455475 699839
rect 455417 699799 455475 699805
rect 8110 699728 8116 699780
rect 8168 699768 8174 699780
rect 422389 699771 422447 699777
rect 422389 699768 422401 699771
rect 8168 699740 422401 699768
rect 8168 699728 8174 699740
rect 422389 699737 422401 699740
rect 422435 699737 422447 699771
rect 433337 699771 433395 699777
rect 433337 699768 433349 699771
rect 422389 699731 422447 699737
rect 431926 699740 433349 699768
rect 14550 699660 14556 699712
rect 14608 699700 14614 699712
rect 431926 699700 431954 699740
rect 433337 699737 433349 699740
rect 433383 699737 433395 699771
rect 433337 699731 433395 699737
rect 14608 699672 431954 699700
rect 14608 699660 14614 699672
rect 3050 671984 3056 672036
rect 3108 672024 3114 672036
rect 35158 672024 35164 672036
rect 3108 671996 35164 672024
rect 3108 671984 3114 671996
rect 35158 671984 35164 671996
rect 35216 671984 35222 672036
rect 3510 658180 3516 658232
rect 3568 658220 3574 658232
rect 14550 658220 14556 658232
rect 3568 658192 14556 658220
rect 3568 658180 3574 658192
rect 14550 658180 14556 658192
rect 14608 658180 14614 658232
rect 3326 619556 3332 619608
rect 3384 619596 3390 619608
rect 161566 619596 161572 619608
rect 3384 619568 161572 619596
rect 3384 619556 3390 619568
rect 161566 619556 161572 619568
rect 161624 619556 161630 619608
rect 3234 607112 3240 607164
rect 3292 607152 3298 607164
rect 40678 607152 40684 607164
rect 3292 607124 40684 607152
rect 3292 607112 3298 607124
rect 40678 607112 40684 607124
rect 40736 607112 40742 607164
rect 3510 567128 3516 567180
rect 3568 567168 3574 567180
rect 161658 567168 161664 567180
rect 3568 567140 161664 567168
rect 3568 567128 3574 567140
rect 161658 567128 161664 567140
rect 161716 567128 161722 567180
rect 3510 554684 3516 554736
rect 3568 554724 3574 554736
rect 43438 554724 43444 554736
rect 3568 554696 43444 554724
rect 3568 554684 3574 554696
rect 43438 554684 43444 554696
rect 43496 554684 43502 554736
rect 3510 516060 3516 516112
rect 3568 516100 3574 516112
rect 161750 516100 161756 516112
rect 3568 516072 161756 516100
rect 3568 516060 3574 516072
rect 161750 516060 161756 516072
rect 161808 516060 161814 516112
rect 3510 502256 3516 502308
rect 3568 502296 3574 502308
rect 14458 502296 14464 502308
rect 3568 502268 14464 502296
rect 3568 502256 3574 502268
rect 14458 502256 14464 502268
rect 14516 502256 14522 502308
rect 3234 463632 3240 463684
rect 3292 463672 3298 463684
rect 32398 463672 32404 463684
rect 3292 463644 32404 463672
rect 3292 463632 3298 463644
rect 32398 463632 32404 463644
rect 32456 463632 32462 463684
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 17218 449868 17224 449880
rect 3384 449840 17224 449868
rect 3384 449828 3390 449840
rect 17218 449828 17224 449840
rect 17276 449828 17282 449880
rect 3510 423580 3516 423632
rect 3568 423620 3574 423632
rect 161842 423620 161848 423632
rect 3568 423592 161848 423620
rect 3568 423580 3574 423592
rect 161842 423580 161848 423592
rect 161900 423580 161906 423632
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 161934 411244 161940 411256
rect 3016 411216 161940 411244
rect 3016 411204 3022 411216
rect 161934 411204 161940 411216
rect 161992 411204 161998 411256
rect 3234 398760 3240 398812
rect 3292 398800 3298 398812
rect 18598 398800 18604 398812
rect 3292 398772 18604 398800
rect 3292 398760 3298 398772
rect 18598 398760 18604 398772
rect 18656 398760 18662 398812
rect 3510 372512 3516 372564
rect 3568 372552 3574 372564
rect 162026 372552 162032 372564
rect 3568 372524 162032 372552
rect 3568 372512 3574 372524
rect 162026 372512 162032 372524
rect 162084 372512 162090 372564
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 79318 346372 79324 346384
rect 3200 346344 79324 346372
rect 3200 346332 3206 346344
rect 79318 346332 79324 346344
rect 79376 346332 79382 346384
rect 3418 306280 3424 306332
rect 3476 306320 3482 306332
rect 29638 306320 29644 306332
rect 3476 306292 29644 306320
rect 3476 306280 3482 306292
rect 29638 306280 29644 306292
rect 29696 306280 29702 306332
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 105538 293944 105544 293956
rect 3108 293916 105544 293944
rect 3108 293904 3114 293916
rect 105538 293904 105544 293916
rect 105596 293904 105602 293956
rect 162302 282276 162308 282328
rect 162360 282316 162366 282328
rect 580258 282316 580264 282328
rect 162360 282288 580264 282316
rect 162360 282276 162366 282288
rect 580258 282276 580264 282288
rect 580316 282276 580322 282328
rect 162118 282208 162124 282260
rect 162176 282248 162182 282260
rect 580350 282248 580356 282260
rect 162176 282220 580356 282248
rect 162176 282208 162182 282220
rect 580350 282208 580356 282220
rect 580408 282208 580414 282260
rect 162210 282140 162216 282192
rect 162268 282180 162274 282192
rect 580442 282180 580448 282192
rect 162268 282152 580448 282180
rect 162268 282140 162274 282152
rect 580442 282140 580448 282152
rect 580500 282140 580506 282192
rect 97258 280100 97264 280152
rect 97316 280140 97322 280152
rect 226702 280140 226708 280152
rect 97316 280112 226708 280140
rect 97316 280100 97322 280112
rect 226702 280100 226708 280112
rect 226760 280100 226766 280152
rect 226978 280100 226984 280152
rect 227036 280140 227042 280152
rect 246298 280140 246304 280152
rect 227036 280112 246304 280140
rect 227036 280100 227042 280112
rect 246298 280100 246304 280112
rect 246356 280100 246362 280152
rect 320082 280100 320088 280152
rect 320140 280140 320146 280152
rect 324041 280143 324099 280149
rect 324041 280140 324053 280143
rect 320140 280112 324053 280140
rect 320140 280100 320146 280112
rect 324041 280109 324053 280112
rect 324087 280109 324099 280143
rect 324041 280103 324099 280109
rect 324133 280143 324191 280149
rect 324133 280109 324145 280143
rect 324179 280140 324191 280143
rect 351914 280140 351920 280152
rect 324179 280112 351920 280140
rect 324179 280109 324191 280112
rect 324133 280103 324191 280109
rect 351914 280100 351920 280112
rect 351972 280100 351978 280152
rect 352558 280100 352564 280152
rect 352616 280140 352622 280152
rect 414934 280140 414940 280152
rect 352616 280112 414940 280140
rect 352616 280100 352622 280112
rect 414934 280100 414940 280112
rect 414992 280100 414998 280152
rect 419442 280100 419448 280152
rect 419500 280140 419506 280152
rect 464338 280140 464344 280152
rect 419500 280112 464344 280140
rect 419500 280100 419506 280112
rect 464338 280100 464344 280112
rect 464396 280100 464402 280152
rect 471882 280100 471888 280152
rect 471940 280140 471946 280152
rect 501874 280140 501880 280152
rect 471940 280112 501880 280140
rect 471940 280100 471946 280112
rect 501874 280100 501880 280112
rect 501932 280100 501938 280152
rect 503622 280100 503628 280152
rect 503680 280140 503686 280152
rect 524874 280140 524880 280152
rect 503680 280112 524880 280140
rect 503680 280100 503686 280112
rect 524874 280100 524880 280112
rect 524932 280100 524938 280152
rect 525150 280100 525156 280152
rect 525208 280140 525214 280152
rect 540238 280140 540244 280152
rect 525208 280112 540244 280140
rect 525208 280100 525214 280112
rect 540238 280100 540244 280112
rect 540296 280100 540302 280152
rect 576854 280100 576860 280152
rect 576912 280140 576918 280152
rect 577682 280140 577688 280152
rect 576912 280112 577688 280140
rect 576912 280100 576918 280112
rect 577682 280100 577688 280112
rect 577740 280100 577746 280152
rect 111702 280032 111708 280084
rect 111760 280072 111766 280084
rect 242066 280072 242072 280084
rect 111760 280044 242072 280072
rect 111760 280032 111766 280044
rect 242066 280032 242072 280044
rect 242124 280032 242130 280084
rect 255406 280032 255412 280084
rect 255464 280072 255470 280084
rect 261662 280072 261668 280084
rect 255464 280044 261668 280072
rect 255464 280032 255470 280044
rect 261662 280032 261668 280044
rect 261720 280032 261726 280084
rect 302878 280032 302884 280084
rect 302936 280072 302942 280084
rect 367278 280072 367284 280084
rect 302936 280044 367284 280072
rect 302936 280032 302942 280044
rect 367278 280032 367284 280044
rect 367336 280032 367342 280084
rect 369762 280032 369768 280084
rect 369820 280072 369826 280084
rect 428642 280072 428648 280084
rect 369820 280044 428648 280072
rect 369820 280032 369826 280044
rect 428642 280032 428648 280044
rect 428700 280032 428706 280084
rect 430482 280032 430488 280084
rect 430540 280072 430546 280084
rect 472066 280072 472072 280084
rect 430540 280044 472072 280072
rect 430540 280032 430546 280044
rect 472066 280032 472072 280044
rect 472124 280032 472130 280084
rect 472618 280032 472624 280084
rect 472676 280072 472682 280084
rect 484854 280072 484860 280084
rect 472676 280044 484860 280072
rect 472676 280032 472682 280044
rect 484854 280032 484860 280044
rect 484912 280032 484918 280084
rect 485682 280032 485688 280084
rect 485740 280072 485746 280084
rect 512086 280072 512092 280084
rect 485740 280044 512092 280072
rect 485740 280032 485746 280044
rect 512086 280032 512092 280044
rect 512144 280032 512150 280084
rect 513282 280032 513288 280084
rect 513340 280072 513346 280084
rect 531682 280072 531688 280084
rect 513340 280044 531688 280072
rect 513340 280032 513346 280044
rect 531682 280032 531688 280044
rect 531740 280032 531746 280084
rect 533430 280032 533436 280084
rect 533488 280072 533494 280084
rect 545298 280072 545304 280084
rect 533488 280044 545304 280072
rect 533488 280032 533494 280044
rect 545298 280032 545304 280044
rect 545356 280032 545362 280084
rect 101398 279964 101404 280016
rect 101456 280004 101462 280016
rect 231854 280004 231860 280016
rect 101456 279976 231860 280004
rect 101456 279964 101462 279976
rect 231854 279964 231860 279976
rect 231912 279964 231918 280016
rect 295978 279964 295984 280016
rect 296036 280004 296042 280016
rect 313550 280004 313556 280016
rect 296036 279976 313556 280004
rect 296036 279964 296042 279976
rect 313550 279964 313556 279976
rect 313608 279964 313614 280016
rect 317417 280007 317475 280013
rect 317417 279973 317429 280007
rect 317463 280004 317475 280007
rect 323854 280004 323860 280016
rect 317463 279976 323860 280004
rect 317463 279973 317475 279976
rect 317417 279967 317475 279973
rect 323854 279964 323860 279976
rect 323912 279964 323918 280016
rect 325697 280007 325755 280013
rect 325697 280004 325709 280007
rect 323964 279976 325709 280004
rect 35158 279896 35164 279948
rect 35216 279936 35222 279948
rect 179874 279936 179880 279948
rect 35216 279908 179880 279936
rect 35216 279896 35222 279908
rect 179874 279896 179880 279908
rect 179932 279896 179938 279948
rect 222838 279896 222844 279948
rect 222896 279936 222902 279948
rect 248874 279936 248880 279948
rect 222896 279908 248880 279936
rect 222896 279896 222902 279908
rect 248874 279896 248880 279908
rect 248932 279896 248938 279948
rect 249058 279896 249064 279948
rect 249116 279936 249122 279948
rect 260834 279936 260840 279948
rect 249116 279908 260840 279936
rect 249116 279896 249122 279908
rect 260834 279896 260840 279908
rect 260892 279896 260898 279948
rect 276658 279896 276664 279948
rect 276716 279936 276722 279948
rect 318794 279936 318800 279948
rect 276716 279908 318800 279936
rect 276716 279896 276722 279908
rect 318794 279896 318800 279908
rect 318852 279896 318858 279948
rect 322198 279896 322204 279948
rect 322256 279936 322262 279948
rect 323964 279936 323992 279976
rect 325697 279973 325709 279976
rect 325743 279973 325755 280007
rect 325697 279967 325755 279973
rect 325786 279964 325792 280016
rect 325844 280004 325850 280016
rect 326338 280004 326344 280016
rect 325844 279976 326344 280004
rect 325844 279964 325850 279976
rect 326338 279964 326344 279976
rect 326396 279964 326402 280016
rect 326433 280007 326491 280013
rect 326433 279973 326445 280007
rect 326479 280004 326491 280007
rect 328914 280004 328920 280016
rect 326479 279976 328920 280004
rect 326479 279973 326491 279976
rect 326433 279967 326491 279973
rect 328914 279964 328920 279976
rect 328972 279964 328978 280016
rect 329098 279964 329104 280016
rect 329156 280004 329162 280016
rect 397914 280004 397920 280016
rect 329156 279976 397920 280004
rect 329156 279964 329162 279976
rect 397914 279964 397920 279976
rect 397972 279964 397978 280016
rect 399478 279964 399484 280016
rect 399536 280004 399542 280016
rect 449066 280004 449072 280016
rect 399536 279976 449072 280004
rect 399536 279964 399542 279976
rect 449066 279964 449072 279976
rect 449124 279964 449130 280016
rect 449802 279964 449808 280016
rect 449860 280004 449866 280016
rect 486510 280004 486516 280016
rect 449860 279976 486516 280004
rect 449860 279964 449866 279976
rect 486510 279964 486516 279976
rect 486568 279964 486574 280016
rect 496722 279964 496728 280016
rect 496780 280004 496786 280016
rect 519722 280004 519728 280016
rect 496780 279976 519728 280004
rect 496780 279964 496786 279976
rect 519722 279964 519728 279976
rect 519780 279964 519786 280016
rect 519817 280007 519875 280013
rect 519817 279973 519829 280007
rect 519863 280004 519875 280007
rect 527450 280004 527456 280016
rect 519863 279976 527456 280004
rect 519863 279973 519875 279976
rect 519817 279967 519875 279973
rect 527450 279964 527456 279976
rect 527508 279964 527514 280016
rect 527545 280007 527603 280013
rect 527545 279973 527557 280007
rect 527591 280004 527603 280007
rect 537662 280004 537668 280016
rect 527591 279976 537668 280004
rect 527591 279973 527603 279976
rect 527545 279967 527603 279973
rect 537662 279964 537668 279976
rect 537720 279964 537726 280016
rect 538122 279964 538128 280016
rect 538180 280004 538186 280016
rect 549530 280004 549536 280016
rect 538180 279976 549536 280004
rect 538180 279964 538186 279976
rect 549530 279964 549536 279976
rect 549588 279964 549594 280016
rect 322256 279908 323992 279936
rect 324041 279939 324099 279945
rect 322256 279896 322262 279908
rect 324041 279905 324053 279939
rect 324087 279936 324099 279939
rect 392854 279936 392860 279948
rect 324087 279908 392860 279936
rect 324087 279905 324099 279908
rect 324041 279899 324099 279905
rect 392854 279896 392860 279908
rect 392912 279896 392918 279948
rect 393958 279896 393964 279948
rect 394016 279936 394022 279948
rect 394016 279908 395476 279936
rect 394016 279896 394022 279908
rect 50338 279828 50344 279880
rect 50396 279868 50402 279880
rect 196066 279868 196072 279880
rect 50396 279840 196072 279868
rect 50396 279828 50402 279840
rect 196066 279828 196072 279840
rect 196124 279828 196130 279880
rect 196618 279828 196624 279880
rect 196676 279868 196682 279880
rect 216674 279868 216680 279880
rect 196676 279840 216680 279868
rect 196676 279828 196682 279840
rect 216674 279828 216680 279840
rect 216732 279828 216738 279880
rect 221458 279828 221464 279880
rect 221516 279868 221522 279880
rect 221516 279840 221688 279868
rect 221516 279828 221522 279840
rect 43438 279760 43444 279812
rect 43496 279800 43502 279812
rect 190914 279800 190920 279812
rect 43496 279772 190920 279800
rect 43496 279760 43502 279772
rect 190914 279760 190920 279772
rect 190972 279760 190978 279812
rect 199378 279760 199384 279812
rect 199436 279800 199442 279812
rect 221550 279800 221556 279812
rect 199436 279772 221556 279800
rect 199436 279760 199442 279772
rect 221550 279760 221556 279772
rect 221608 279760 221614 279812
rect 221660 279800 221688 279840
rect 221734 279828 221740 279880
rect 221792 279868 221798 279880
rect 249794 279868 249800 279880
rect 221792 279840 249800 279868
rect 221792 279828 221798 279840
rect 249794 279828 249800 279840
rect 249852 279828 249858 279880
rect 252002 279828 252008 279880
rect 252060 279868 252066 279880
rect 278774 279868 278780 279880
rect 252060 279840 278780 279868
rect 252060 279828 252066 279840
rect 278774 279828 278780 279840
rect 278832 279828 278838 279880
rect 309134 279828 309140 279880
rect 309192 279868 309198 279880
rect 310146 279868 310152 279880
rect 309192 279840 310152 279868
rect 309192 279828 309198 279840
rect 310146 279828 310152 279840
rect 310204 279828 310210 279880
rect 313182 279828 313188 279880
rect 313240 279868 313246 279880
rect 387794 279868 387800 279880
rect 313240 279840 387800 279868
rect 313240 279828 313246 279840
rect 387794 279828 387800 279840
rect 387852 279828 387858 279880
rect 387904 279840 393314 279868
rect 244550 279800 244556 279812
rect 221660 279772 244556 279800
rect 244550 279760 244556 279772
rect 244608 279760 244614 279812
rect 244918 279760 244924 279812
rect 244976 279800 244982 279812
rect 283742 279800 283748 279812
rect 244976 279772 283748 279800
rect 244976 279760 244982 279772
rect 283742 279760 283748 279772
rect 283800 279760 283806 279812
rect 306282 279760 306288 279812
rect 306340 279800 306346 279812
rect 382550 279800 382556 279812
rect 306340 279772 382556 279800
rect 306340 279760 306346 279772
rect 382550 279760 382556 279772
rect 382608 279760 382614 279812
rect 384390 279760 384396 279812
rect 384448 279800 384454 279812
rect 387904 279800 387932 279840
rect 384448 279772 387932 279800
rect 384448 279760 384454 279772
rect 389818 279760 389824 279812
rect 389876 279800 389882 279812
rect 390554 279800 390560 279812
rect 389876 279772 390560 279800
rect 389876 279760 389882 279772
rect 390554 279760 390560 279772
rect 390612 279760 390618 279812
rect 393286 279800 393314 279840
rect 394694 279828 394700 279880
rect 394752 279868 394758 279880
rect 395338 279868 395344 279880
rect 394752 279840 395344 279868
rect 394752 279828 394758 279840
rect 395338 279828 395344 279840
rect 395396 279828 395402 279880
rect 395448 279868 395476 279908
rect 400122 279896 400128 279948
rect 400180 279936 400186 279948
rect 450722 279936 450728 279948
rect 400180 279908 450728 279936
rect 400180 279896 400186 279908
rect 450722 279896 450728 279908
rect 450780 279896 450786 279948
rect 454678 279896 454684 279948
rect 454736 279936 454742 279948
rect 463694 279936 463700 279948
rect 454736 279908 463700 279936
rect 454736 279896 454742 279908
rect 463694 279896 463700 279908
rect 463752 279896 463758 279948
rect 466362 279896 466368 279948
rect 466420 279936 466426 279948
rect 497642 279936 497648 279948
rect 466420 279908 497648 279936
rect 466420 279896 466426 279908
rect 497642 279896 497648 279908
rect 497700 279896 497706 279948
rect 502242 279896 502248 279948
rect 502300 279936 502306 279948
rect 524046 279936 524052 279948
rect 502300 279908 524052 279936
rect 502300 279896 502306 279908
rect 524046 279896 524052 279908
rect 524104 279896 524110 279948
rect 525058 279896 525064 279948
rect 525116 279936 525122 279948
rect 539594 279936 539600 279948
rect 525116 279908 539600 279936
rect 525116 279896 525122 279908
rect 539594 279896 539600 279908
rect 539652 279896 539658 279948
rect 542998 279896 543004 279948
rect 543056 279936 543062 279948
rect 552934 279936 552940 279948
rect 543056 279908 552940 279936
rect 543056 279896 543062 279908
rect 552934 279896 552940 279908
rect 552992 279896 552998 279948
rect 445754 279868 445760 279880
rect 395448 279840 445760 279868
rect 445754 279828 445760 279840
rect 445812 279828 445818 279880
rect 451182 279828 451188 279880
rect 451240 279868 451246 279880
rect 487338 279868 487344 279880
rect 451240 279840 487344 279868
rect 451240 279828 451246 279840
rect 487338 279828 487344 279840
rect 487396 279828 487402 279880
rect 489822 279828 489828 279880
rect 489880 279868 489886 279880
rect 514754 279868 514760 279880
rect 489880 279840 514760 279868
rect 489880 279828 489886 279840
rect 514754 279828 514760 279840
rect 514812 279828 514818 279880
rect 516042 279828 516048 279880
rect 516100 279868 516106 279880
rect 534258 279868 534264 279880
rect 516100 279840 534264 279868
rect 516100 279828 516106 279840
rect 534258 279828 534264 279840
rect 534316 279828 534322 279880
rect 536742 279828 536748 279880
rect 536800 279868 536806 279880
rect 548702 279868 548708 279880
rect 536800 279840 548708 279868
rect 536800 279828 536806 279840
rect 548702 279828 548708 279840
rect 548760 279828 548766 279880
rect 438854 279800 438860 279812
rect 393286 279772 438860 279800
rect 438854 279760 438860 279772
rect 438912 279760 438918 279812
rect 440142 279760 440148 279812
rect 440200 279800 440206 279812
rect 478874 279800 478880 279812
rect 440200 279772 478880 279800
rect 440200 279760 440206 279772
rect 478874 279760 478880 279772
rect 478932 279760 478938 279812
rect 482922 279760 482928 279812
rect 482980 279800 482986 279812
rect 509510 279800 509516 279812
rect 482980 279772 509516 279800
rect 482980 279760 482986 279772
rect 509510 279760 509516 279772
rect 509568 279760 509574 279812
rect 514662 279760 514668 279812
rect 514720 279800 514726 279812
rect 532694 279800 532700 279812
rect 514720 279772 532700 279800
rect 514720 279760 514726 279772
rect 532694 279760 532700 279772
rect 532752 279760 532758 279812
rect 533338 279760 533344 279812
rect 533396 279800 533402 279812
rect 546126 279800 546132 279812
rect 533396 279772 546132 279800
rect 533396 279760 533402 279772
rect 546126 279760 546132 279772
rect 546184 279760 546190 279812
rect 547138 279760 547144 279812
rect 547196 279800 547202 279812
rect 555510 279800 555516 279812
rect 547196 279772 555516 279800
rect 547196 279760 547202 279772
rect 555510 279760 555516 279772
rect 555568 279760 555574 279812
rect 36538 279692 36544 279744
rect 36596 279732 36602 279744
rect 185854 279732 185860 279744
rect 36596 279704 185860 279732
rect 36596 279692 36602 279704
rect 185854 279692 185860 279704
rect 185912 279692 185918 279744
rect 208486 279692 208492 279744
rect 208544 279732 208550 279744
rect 251450 279732 251456 279744
rect 208544 279704 251456 279732
rect 208544 279692 208550 279704
rect 251450 279692 251456 279704
rect 251508 279692 251514 279744
rect 251818 279692 251824 279744
rect 251876 279732 251882 279744
rect 254854 279732 254860 279744
rect 251876 279704 254860 279732
rect 251876 279692 251882 279704
rect 254854 279692 254860 279704
rect 254912 279692 254918 279744
rect 254949 279735 255007 279741
rect 254949 279701 254961 279735
rect 254995 279732 255007 279735
rect 281534 279732 281540 279744
rect 254995 279704 281540 279732
rect 254995 279701 255007 279704
rect 254949 279695 255007 279701
rect 281534 279692 281540 279704
rect 281592 279692 281598 279744
rect 299382 279692 299388 279744
rect 299440 279732 299446 279744
rect 377490 279732 377496 279744
rect 299440 279704 377496 279732
rect 299440 279692 299446 279704
rect 377490 279692 377496 279704
rect 377548 279692 377554 279744
rect 377582 279692 377588 279744
rect 377640 279732 377646 279744
rect 433702 279732 433708 279744
rect 377640 279704 433708 279732
rect 377640 279692 377646 279704
rect 433702 279692 433708 279704
rect 433760 279692 433766 279744
rect 437382 279692 437388 279744
rect 437440 279732 437446 279744
rect 477126 279732 477132 279744
rect 437440 279704 477132 279732
rect 437440 279692 437446 279704
rect 477126 279692 477132 279704
rect 477184 279692 477190 279744
rect 479518 279692 479524 279744
rect 479576 279732 479582 279744
rect 506934 279732 506940 279744
rect 479576 279704 506940 279732
rect 479576 279692 479582 279704
rect 506934 279692 506940 279704
rect 506992 279692 506998 279744
rect 507762 279692 507768 279744
rect 507820 279732 507826 279744
rect 519449 279735 519507 279741
rect 519449 279732 519461 279735
rect 507820 279704 519461 279732
rect 507820 279692 507826 279704
rect 519449 279701 519461 279704
rect 519495 279701 519507 279735
rect 519449 279695 519507 279701
rect 519538 279692 519544 279744
rect 519596 279732 519602 279744
rect 526530 279732 526536 279744
rect 519596 279704 526536 279732
rect 519596 279692 519602 279704
rect 526530 279692 526536 279704
rect 526588 279692 526594 279744
rect 535362 279692 535368 279744
rect 535420 279732 535426 279744
rect 548058 279732 548064 279744
rect 535420 279704 548064 279732
rect 535420 279692 535426 279704
rect 548058 279692 548064 279704
rect 548116 279692 548122 279744
rect 549162 279692 549168 279744
rect 549220 279732 549226 279744
rect 558086 279732 558092 279744
rect 549220 279704 558092 279732
rect 549220 279692 549226 279704
rect 558086 279692 558092 279704
rect 558144 279692 558150 279744
rect 29638 279624 29644 279676
rect 29696 279664 29702 279676
rect 180886 279664 180892 279676
rect 29696 279636 180892 279664
rect 29696 279624 29702 279636
rect 180886 279624 180892 279636
rect 180944 279624 180950 279676
rect 187694 279624 187700 279676
rect 187752 279664 187758 279676
rect 188338 279664 188344 279676
rect 187752 279636 188344 279664
rect 187752 279624 187758 279636
rect 188338 279624 188344 279636
rect 188396 279624 188402 279676
rect 200758 279624 200764 279676
rect 200816 279664 200822 279676
rect 224126 279664 224132 279676
rect 200816 279636 224132 279664
rect 200816 279624 200822 279636
rect 224126 279624 224132 279636
rect 224184 279624 224190 279676
rect 233878 279624 233884 279676
rect 233936 279664 233942 279676
rect 286318 279664 286324 279676
rect 233936 279636 286324 279664
rect 233936 279624 233942 279636
rect 286318 279624 286324 279636
rect 286376 279624 286382 279676
rect 293218 279624 293224 279676
rect 293276 279664 293282 279676
rect 372614 279664 372620 279676
rect 293276 279636 372620 279664
rect 293276 279624 293282 279636
rect 372614 279624 372620 279636
rect 372672 279624 372678 279676
rect 373258 279624 373264 279676
rect 373316 279664 373322 279676
rect 425609 279667 425667 279673
rect 425609 279664 425621 279667
rect 373316 279636 425621 279664
rect 373316 279624 373322 279636
rect 425609 279633 425621 279636
rect 425655 279633 425667 279667
rect 425609 279627 425667 279633
rect 425698 279624 425704 279676
rect 425756 279664 425762 279676
rect 431126 279664 431132 279676
rect 425756 279636 431132 279664
rect 425756 279624 425762 279636
rect 431126 279624 431132 279636
rect 431184 279624 431190 279676
rect 433242 279624 433248 279676
rect 433300 279664 433306 279676
rect 473722 279664 473728 279676
rect 433300 279636 473728 279664
rect 433300 279624 433306 279636
rect 473722 279624 473728 279636
rect 473780 279624 473786 279676
rect 480898 279624 480904 279676
rect 480956 279664 480962 279676
rect 507854 279664 507860 279676
rect 480956 279636 507860 279664
rect 480956 279624 480962 279636
rect 507854 279624 507860 279636
rect 507912 279624 507918 279676
rect 509142 279624 509148 279676
rect 509200 279664 509206 279676
rect 529106 279664 529112 279676
rect 509200 279636 529112 279664
rect 509200 279624 509206 279636
rect 529106 279624 529112 279636
rect 529164 279624 529170 279676
rect 529842 279624 529848 279676
rect 529900 279664 529906 279676
rect 543734 279664 543740 279676
rect 529900 279636 543740 279664
rect 529900 279624 529906 279636
rect 543734 279624 543740 279636
rect 543792 279624 543798 279676
rect 544378 279624 544384 279676
rect 544436 279664 544442 279676
rect 553854 279664 553860 279676
rect 544436 279636 553860 279664
rect 544436 279624 544442 279636
rect 553854 279624 553860 279636
rect 553912 279624 553918 279676
rect 558178 279624 558184 279676
rect 558236 279664 558242 279676
rect 562318 279664 562324 279676
rect 558236 279636 562324 279664
rect 558236 279624 558242 279636
rect 562318 279624 562324 279636
rect 562376 279624 562382 279676
rect 572714 279624 572720 279676
rect 572772 279664 572778 279676
rect 573450 279664 573456 279676
rect 572772 279636 573456 279664
rect 572772 279624 572778 279636
rect 573450 279624 573456 279636
rect 573508 279624 573514 279676
rect 582282 279624 582288 279676
rect 582340 279664 582346 279676
rect 583021 279667 583079 279673
rect 583021 279664 583033 279667
rect 582340 279636 583033 279664
rect 582340 279624 582346 279636
rect 583021 279633 583033 279636
rect 583067 279633 583079 279667
rect 583021 279627 583079 279633
rect 18598 279556 18604 279608
rect 18656 279596 18662 279608
rect 173066 279596 173072 279608
rect 18656 279568 173072 279596
rect 18656 279556 18662 279568
rect 173066 279556 173072 279568
rect 173124 279556 173130 279608
rect 195238 279556 195244 279608
rect 195296 279596 195302 279608
rect 211338 279596 211344 279608
rect 195296 279568 211344 279596
rect 195296 279556 195302 279568
rect 211338 279556 211344 279568
rect 211396 279556 211402 279608
rect 214558 279556 214564 279608
rect 214616 279596 214622 279608
rect 239490 279596 239496 279608
rect 214616 279568 239496 279596
rect 214616 279556 214622 279568
rect 239490 279556 239496 279568
rect 239548 279556 239554 279608
rect 242802 279556 242808 279608
rect 242860 279596 242866 279608
rect 317417 279599 317475 279605
rect 317417 279596 317429 279599
rect 242860 279568 317429 279596
rect 242860 279556 242866 279568
rect 317417 279565 317429 279568
rect 317463 279565 317475 279599
rect 317417 279559 317475 279565
rect 317506 279556 317512 279608
rect 317564 279596 317570 279608
rect 321554 279596 321560 279608
rect 317564 279568 321560 279596
rect 317564 279556 317570 279568
rect 321554 279556 321560 279568
rect 321612 279556 321618 279608
rect 327074 279556 327080 279608
rect 327132 279596 327138 279608
rect 328086 279596 328092 279608
rect 327132 279568 328092 279596
rect 327132 279556 327138 279568
rect 328086 279556 328092 279568
rect 328144 279556 328150 279608
rect 334066 279556 334072 279608
rect 334124 279596 334130 279608
rect 334894 279596 334900 279608
rect 334124 279568 334900 279596
rect 334124 279556 334130 279568
rect 334894 279556 334900 279568
rect 334952 279556 334958 279608
rect 334989 279599 335047 279605
rect 334989 279565 335001 279599
rect 335035 279596 335047 279599
rect 403158 279596 403164 279608
rect 335035 279568 403164 279596
rect 335035 279565 335047 279568
rect 334989 279559 335047 279565
rect 403158 279556 403164 279568
rect 403216 279556 403222 279608
rect 407758 279556 407764 279608
rect 407816 279596 407822 279608
rect 410702 279596 410708 279608
rect 407816 279568 410708 279596
rect 407816 279556 407822 279568
rect 410702 279556 410708 279568
rect 410760 279556 410766 279608
rect 410797 279599 410855 279605
rect 410797 279565 410809 279599
rect 410843 279596 410855 279599
rect 454126 279596 454132 279608
rect 410843 279568 454132 279596
rect 410843 279565 410855 279568
rect 410797 279559 410855 279565
rect 454126 279556 454132 279568
rect 454184 279556 454190 279608
rect 458082 279556 458088 279608
rect 458140 279596 458146 279608
rect 492674 279596 492680 279608
rect 458140 279568 492680 279596
rect 458140 279556 458146 279568
rect 492674 279556 492680 279568
rect 492732 279556 492738 279608
rect 493318 279556 493324 279608
rect 493376 279596 493382 279608
rect 517514 279596 517520 279608
rect 493376 279568 517520 279596
rect 493376 279556 493382 279568
rect 517514 279556 517520 279568
rect 517572 279556 517578 279608
rect 522942 279556 522948 279608
rect 523000 279596 523006 279608
rect 538490 279596 538496 279608
rect 523000 279568 538496 279596
rect 523000 279556 523006 279568
rect 538490 279556 538496 279568
rect 538548 279556 538554 279608
rect 539502 279556 539508 279608
rect 539560 279596 539566 279608
rect 550634 279596 550640 279608
rect 539560 279568 550640 279596
rect 539560 279556 539566 279568
rect 550634 279556 550640 279568
rect 550692 279556 550698 279608
rect 558270 279556 558276 279608
rect 558328 279596 558334 279608
rect 563238 279596 563244 279608
rect 558328 279568 563244 279596
rect 558328 279556 558334 279568
rect 563238 279556 563244 279568
rect 563296 279556 563302 279608
rect 572622 279556 572628 279608
rect 572680 279596 572686 279608
rect 574278 279596 574284 279608
rect 572680 279568 574284 279596
rect 572680 279556 572686 279568
rect 574278 279556 574284 279568
rect 574336 279556 574342 279608
rect 17218 279488 17224 279540
rect 17276 279528 17282 279540
rect 173894 279528 173900 279540
rect 17276 279500 173900 279528
rect 17276 279488 17282 279500
rect 173894 279488 173900 279500
rect 173952 279488 173958 279540
rect 191098 279488 191104 279540
rect 191156 279528 191162 279540
rect 201126 279528 201132 279540
rect 191156 279500 201132 279528
rect 191156 279488 191162 279500
rect 201126 279488 201132 279500
rect 201184 279488 201190 279540
rect 203518 279488 203524 279540
rect 203576 279528 203582 279540
rect 229370 279528 229376 279540
rect 203576 279500 229376 279528
rect 203576 279488 203582 279500
rect 229370 279488 229376 279500
rect 229428 279488 229434 279540
rect 251910 279488 251916 279540
rect 251968 279528 251974 279540
rect 254949 279531 255007 279537
rect 254949 279528 254961 279531
rect 251968 279500 254961 279528
rect 251968 279488 251974 279500
rect 254949 279497 254961 279500
rect 254995 279497 255007 279531
rect 254949 279491 255007 279497
rect 255041 279531 255099 279537
rect 255041 279497 255053 279531
rect 255087 279528 255099 279531
rect 341702 279528 341708 279540
rect 255087 279500 341708 279528
rect 255087 279497 255099 279500
rect 255041 279491 255099 279497
rect 341702 279488 341708 279500
rect 341760 279488 341766 279540
rect 342898 279488 342904 279540
rect 342956 279528 342962 279540
rect 344278 279528 344284 279540
rect 342956 279500 344284 279528
rect 342956 279488 342962 279500
rect 344278 279488 344284 279500
rect 344336 279488 344342 279540
rect 349062 279488 349068 279540
rect 349120 279528 349126 279540
rect 413278 279528 413284 279540
rect 349120 279500 413284 279528
rect 349120 279488 349126 279500
rect 413278 279488 413284 279500
rect 413336 279488 413342 279540
rect 415302 279488 415308 279540
rect 415360 279528 415366 279540
rect 461026 279528 461032 279540
rect 415360 279500 461032 279528
rect 415360 279488 415366 279500
rect 461026 279488 461032 279500
rect 461084 279488 461090 279540
rect 464430 279488 464436 279540
rect 464488 279528 464494 279540
rect 466086 279528 466092 279540
rect 464488 279500 466092 279528
rect 464488 279488 464494 279500
rect 466086 279488 466092 279500
rect 466144 279488 466150 279540
rect 467098 279488 467104 279540
rect 467156 279528 467162 279540
rect 469490 279528 469496 279540
rect 467156 279500 469496 279528
rect 467156 279488 467162 279500
rect 469490 279488 469496 279500
rect 469548 279488 469554 279540
rect 469585 279531 469643 279537
rect 469585 279497 469597 279531
rect 469631 279528 469643 279531
rect 494146 279528 494152 279540
rect 469631 279500 494152 279528
rect 469631 279497 469643 279500
rect 469585 279491 469643 279497
rect 494146 279488 494152 279500
rect 494204 279488 494210 279540
rect 495342 279488 495348 279540
rect 495400 279528 495406 279540
rect 518894 279528 518900 279540
rect 495400 279500 518900 279528
rect 495400 279488 495406 279500
rect 518894 279488 518900 279500
rect 518952 279488 518958 279540
rect 520182 279488 520188 279540
rect 520240 279528 520246 279540
rect 536834 279528 536840 279540
rect 520240 279500 536840 279528
rect 520240 279488 520246 279500
rect 536834 279488 536840 279500
rect 536892 279488 536898 279540
rect 540882 279488 540888 279540
rect 540940 279528 540946 279540
rect 552106 279528 552112 279540
rect 540940 279500 552112 279528
rect 540940 279488 540946 279500
rect 552106 279488 552112 279500
rect 552164 279488 552170 279540
rect 554682 279488 554688 279540
rect 554740 279528 554746 279540
rect 561674 279528 561680 279540
rect 554740 279500 561680 279528
rect 554740 279488 554746 279500
rect 561674 279488 561680 279500
rect 561732 279488 561738 279540
rect 569218 279488 569224 279540
rect 569276 279528 569282 279540
rect 571702 279528 571708 279540
rect 569276 279500 571708 279528
rect 569276 279488 569282 279500
rect 571702 279488 571708 279500
rect 571760 279488 571766 279540
rect 7558 279420 7564 279472
rect 7616 279460 7622 279472
rect 167086 279460 167092 279472
rect 7616 279432 167092 279460
rect 7616 279420 7622 279432
rect 167086 279420 167092 279432
rect 167144 279420 167150 279472
rect 169754 279420 169760 279472
rect 169812 279460 169818 279472
rect 170490 279460 170496 279472
rect 169812 279432 170496 279460
rect 169812 279420 169818 279432
rect 170490 279420 170496 279432
rect 170548 279420 170554 279472
rect 180058 279420 180064 279472
rect 180116 279460 180122 279472
rect 190086 279460 190092 279472
rect 180116 279432 190092 279460
rect 180116 279420 180122 279432
rect 190086 279420 190092 279432
rect 190144 279420 190150 279472
rect 192478 279420 192484 279472
rect 192536 279460 192542 279472
rect 206278 279460 206284 279472
rect 192536 279432 206284 279460
rect 192536 279420 192542 279432
rect 206278 279420 206284 279432
rect 206336 279420 206342 279472
rect 206370 279420 206376 279472
rect 206428 279460 206434 279472
rect 234614 279460 234620 279472
rect 206428 279432 234620 279460
rect 206428 279420 206434 279432
rect 234614 279420 234620 279432
rect 234672 279420 234678 279472
rect 242710 279420 242716 279472
rect 242768 279460 242774 279472
rect 336734 279460 336740 279472
rect 242768 279432 336740 279460
rect 242768 279420 242774 279432
rect 336734 279420 336740 279432
rect 336792 279420 336798 279472
rect 342162 279420 342168 279472
rect 342220 279460 342226 279472
rect 408126 279460 408132 279472
rect 342220 279432 408132 279460
rect 342220 279420 342226 279432
rect 408126 279420 408132 279432
rect 408184 279420 408190 279472
rect 412542 279420 412548 279472
rect 412600 279460 412606 279472
rect 459554 279460 459560 279472
rect 412600 279432 459560 279460
rect 412600 279420 412606 279432
rect 459554 279420 459560 279432
rect 459612 279420 459618 279472
rect 464338 279420 464344 279472
rect 464396 279460 464402 279472
rect 466914 279460 466920 279472
rect 464396 279432 466920 279460
rect 464396 279420 464402 279432
rect 466914 279420 466920 279432
rect 466972 279420 466978 279472
rect 467742 279420 467748 279472
rect 467800 279460 467806 279472
rect 499574 279460 499580 279472
rect 467800 279432 499580 279460
rect 467800 279420 467806 279432
rect 499574 279420 499580 279432
rect 499632 279420 499638 279472
rect 500862 279420 500868 279472
rect 500920 279460 500926 279472
rect 523126 279460 523132 279472
rect 500920 279432 523132 279460
rect 500920 279420 500926 279432
rect 523126 279420 523132 279432
rect 523184 279420 523190 279472
rect 526438 279420 526444 279472
rect 526496 279460 526502 279472
rect 541066 279460 541072 279472
rect 526496 279432 541072 279460
rect 526496 279420 526502 279432
rect 541066 279420 541072 279432
rect 541124 279420 541130 279472
rect 545022 279420 545028 279472
rect 545080 279460 545086 279472
rect 554774 279460 554780 279472
rect 545080 279432 554780 279460
rect 545080 279420 545086 279432
rect 554774 279420 554780 279432
rect 554832 279420 554838 279472
rect 557442 279420 557448 279472
rect 557500 279460 557506 279472
rect 564066 279460 564072 279472
rect 557500 279432 564072 279460
rect 557500 279420 557506 279432
rect 564066 279420 564072 279432
rect 564124 279420 564130 279472
rect 565722 279420 565728 279472
rect 565780 279460 565786 279472
rect 570046 279460 570052 279472
rect 565780 279432 570052 279460
rect 565780 279420 565786 279432
rect 570046 279420 570052 279432
rect 570104 279420 570110 279472
rect 118602 279352 118608 279404
rect 118660 279392 118666 279404
rect 247126 279392 247132 279404
rect 118660 279364 247132 279392
rect 118660 279352 118666 279364
rect 247126 279352 247132 279364
rect 247184 279352 247190 279404
rect 249702 279352 249708 279404
rect 249760 279392 249766 279404
rect 255041 279395 255099 279401
rect 255041 279392 255053 279395
rect 249760 279364 255053 279392
rect 249760 279352 249766 279364
rect 255041 279361 255053 279364
rect 255087 279361 255099 279395
rect 255041 279355 255099 279361
rect 269114 279352 269120 279404
rect 269172 279392 269178 279404
rect 270126 279392 270132 279404
rect 269172 279364 270132 279392
rect 269172 279352 269178 279364
rect 270126 279352 270132 279364
rect 270184 279352 270190 279404
rect 300118 279352 300124 279404
rect 300176 279392 300182 279404
rect 357066 279392 357072 279404
rect 300176 279364 357072 279392
rect 300176 279352 300182 279364
rect 357066 279352 357072 279364
rect 357124 279352 357130 279404
rect 358814 279352 358820 279404
rect 358872 279392 358878 279404
rect 359550 279392 359556 279404
rect 358872 279364 359556 279392
rect 358872 279352 358878 279364
rect 359550 279352 359556 279364
rect 359608 279352 359614 279404
rect 359829 279395 359887 279401
rect 359829 279361 359841 279395
rect 359875 279392 359887 279395
rect 418338 279392 418344 279404
rect 359875 279364 418344 279392
rect 359875 279361 359887 279364
rect 359829 279355 359887 279361
rect 418338 279352 418344 279364
rect 418396 279352 418402 279404
rect 421558 279352 421564 279404
rect 421616 279392 421622 279404
rect 426066 279392 426072 279404
rect 421616 279364 426072 279392
rect 421616 279352 421622 279364
rect 426066 279352 426072 279364
rect 426124 279352 426130 279404
rect 431218 279352 431224 279404
rect 431276 279392 431282 279404
rect 436278 279392 436284 279404
rect 431276 279364 436284 279392
rect 431276 279352 431282 279364
rect 436278 279352 436284 279364
rect 436336 279352 436342 279404
rect 444282 279352 444288 279404
rect 444340 279392 444346 279404
rect 482278 279392 482284 279404
rect 444340 279364 482284 279392
rect 444340 279352 444346 279364
rect 482278 279352 482284 279364
rect 482336 279352 482342 279404
rect 487062 279352 487068 279404
rect 487120 279392 487126 279404
rect 512914 279392 512920 279404
rect 487120 279364 512920 279392
rect 487120 279352 487126 279364
rect 512914 279352 512920 279364
rect 512972 279352 512978 279404
rect 515950 279352 515956 279404
rect 516008 279392 516014 279404
rect 533522 279392 533528 279404
rect 516008 279364 533528 279392
rect 516008 279352 516014 279364
rect 533522 279352 533528 279364
rect 533580 279352 533586 279404
rect 108298 279284 108304 279336
rect 108356 279324 108362 279336
rect 236914 279324 236920 279336
rect 108356 279296 236920 279324
rect 108356 279284 108362 279296
rect 236914 279284 236920 279296
rect 236972 279284 236978 279336
rect 316034 279284 316040 279336
rect 316092 279324 316098 279336
rect 316954 279324 316960 279336
rect 316092 279296 316960 279324
rect 316092 279284 316098 279296
rect 316954 279284 316960 279296
rect 317012 279284 317018 279336
rect 323578 279284 323584 279336
rect 323636 279324 323642 279336
rect 346854 279324 346860 279336
rect 323636 279296 346860 279324
rect 323636 279284 323642 279296
rect 346854 279284 346860 279296
rect 346912 279284 346918 279336
rect 358722 279284 358728 279336
rect 358780 279324 358786 279336
rect 420086 279324 420092 279336
rect 358780 279296 420092 279324
rect 358780 279284 358786 279296
rect 420086 279284 420092 279296
rect 420144 279284 420150 279336
rect 425609 279327 425667 279333
rect 425609 279293 425621 279327
rect 425655 279324 425667 279327
rect 430574 279324 430580 279336
rect 425655 279296 430580 279324
rect 425655 279293 425667 279296
rect 425609 279287 425667 279293
rect 430574 279284 430580 279296
rect 430632 279284 430638 279336
rect 461578 279284 461584 279336
rect 461636 279324 461642 279336
rect 491662 279324 491668 279336
rect 461636 279296 491668 279324
rect 461636 279284 461642 279296
rect 491662 279284 491668 279296
rect 491720 279284 491726 279336
rect 501598 279284 501604 279336
rect 501656 279324 501662 279336
rect 520642 279324 520648 279336
rect 501656 279296 520648 279324
rect 501656 279284 501662 279296
rect 520642 279284 520648 279296
rect 520700 279284 520706 279336
rect 527082 279284 527088 279336
rect 527140 279324 527146 279336
rect 541894 279324 541900 279336
rect 527140 279296 541900 279324
rect 527140 279284 527146 279296
rect 541894 279284 541900 279296
rect 541952 279284 541958 279336
rect 125502 279216 125508 279268
rect 125560 279256 125566 279268
rect 252554 279256 252560 279268
rect 125560 279228 252560 279256
rect 125560 279216 125566 279228
rect 252554 279216 252560 279228
rect 252612 279216 252618 279268
rect 307018 279216 307024 279268
rect 307076 279256 307082 279268
rect 362126 279256 362132 279268
rect 307076 279228 362132 279256
rect 307076 279216 307082 279228
rect 362126 279216 362132 279228
rect 362184 279216 362190 279268
rect 364978 279216 364984 279268
rect 365036 279256 365042 279268
rect 423674 279256 423680 279268
rect 365036 279228 423680 279256
rect 365036 279216 365042 279228
rect 423674 279216 423680 279228
rect 423732 279216 423738 279268
rect 454770 279216 454776 279268
rect 454828 279256 454834 279268
rect 458450 279256 458456 279268
rect 454828 279228 458456 279256
rect 454828 279216 454834 279228
rect 458450 279216 458456 279228
rect 458508 279216 458514 279268
rect 460290 279216 460296 279268
rect 460348 279256 460354 279268
rect 489086 279256 489092 279268
rect 460348 279228 489092 279256
rect 460348 279216 460354 279228
rect 489086 279216 489092 279228
rect 489144 279216 489150 279268
rect 502978 279216 502984 279268
rect 503036 279256 503042 279268
rect 506106 279256 506112 279268
rect 503036 279228 506112 279256
rect 503036 279216 503042 279228
rect 506106 279216 506112 279228
rect 506164 279216 506170 279268
rect 511902 279216 511908 279268
rect 511960 279256 511966 279268
rect 530854 279256 530860 279268
rect 511960 279228 530860 279256
rect 511960 279216 511966 279228
rect 530854 279216 530860 279228
rect 530912 279216 530918 279268
rect 531222 279216 531228 279268
rect 531280 279256 531286 279268
rect 544470 279256 544476 279268
rect 531280 279228 544476 279256
rect 531280 279216 531286 279228
rect 544470 279216 544476 279228
rect 544528 279216 544534 279268
rect 548518 279216 548524 279268
rect 548576 279256 548582 279268
rect 556338 279256 556344 279268
rect 548576 279228 556344 279256
rect 548576 279216 548582 279228
rect 556338 279216 556344 279228
rect 556396 279216 556402 279268
rect 561582 279216 561588 279268
rect 561640 279256 561646 279268
rect 566642 279256 566648 279268
rect 561640 279228 566648 279256
rect 561640 279216 561646 279228
rect 566642 279216 566648 279228
rect 566700 279216 566706 279268
rect 94498 279148 94504 279200
rect 94556 279188 94562 279200
rect 219066 279188 219072 279200
rect 94556 279160 219072 279188
rect 94556 279148 94562 279160
rect 219066 279148 219072 279160
rect 219124 279148 219130 279200
rect 313918 279148 313924 279200
rect 313976 279188 313982 279200
rect 331490 279188 331496 279200
rect 313976 279160 331496 279188
rect 313976 279148 313982 279160
rect 331490 279148 331496 279160
rect 331548 279148 331554 279200
rect 333882 279148 333888 279200
rect 333940 279188 333946 279200
rect 334989 279191 335047 279197
rect 334989 279188 335001 279191
rect 333940 279160 335001 279188
rect 333940 279148 333946 279160
rect 334989 279157 335001 279160
rect 335035 279157 335047 279191
rect 334989 279151 335047 279157
rect 356698 279148 356704 279200
rect 356756 279188 356762 279200
rect 359829 279191 359887 279197
rect 359829 279188 359841 279191
rect 356756 279160 359841 279188
rect 356756 279148 356762 279160
rect 359829 279157 359841 279160
rect 359875 279157 359887 279191
rect 359829 279151 359887 279157
rect 366358 279148 366364 279200
rect 366416 279188 366422 279200
rect 425146 279188 425152 279200
rect 366416 279160 425152 279188
rect 366416 279148 366422 279160
rect 425146 279148 425152 279160
rect 425204 279148 425210 279200
rect 449158 279148 449164 279200
rect 449216 279188 449222 279200
rect 471146 279188 471152 279200
rect 449216 279160 471152 279188
rect 449216 279148 449222 279160
rect 471146 279148 471152 279160
rect 471204 279148 471210 279200
rect 479610 279148 479616 279200
rect 479668 279188 479674 279200
rect 505278 279188 505284 279200
rect 479668 279160 505284 279188
rect 479668 279148 479674 279160
rect 505278 279148 505284 279160
rect 505336 279148 505342 279200
rect 517422 279148 517428 279200
rect 517480 279188 517486 279200
rect 535086 279188 535092 279200
rect 517480 279160 535092 279188
rect 517480 279148 517486 279160
rect 535086 279148 535092 279160
rect 535144 279148 535150 279200
rect 90358 279080 90364 279132
rect 90416 279120 90422 279132
rect 208854 279120 208860 279132
rect 90416 279092 208860 279120
rect 90416 279080 90422 279092
rect 208854 279080 208860 279092
rect 208912 279080 208918 279132
rect 320818 279080 320824 279132
rect 320876 279120 320882 279132
rect 324133 279123 324191 279129
rect 324133 279120 324145 279123
rect 320876 279092 324145 279120
rect 320876 279080 320882 279092
rect 324133 279089 324145 279092
rect 324179 279089 324191 279123
rect 324133 279083 324191 279089
rect 379422 279080 379428 279132
rect 379480 279120 379486 279132
rect 435450 279120 435456 279132
rect 379480 279092 435456 279120
rect 379480 279080 379486 279092
rect 435450 279080 435456 279092
rect 435508 279080 435514 279132
rect 456058 279080 456064 279132
rect 456116 279120 456122 279132
rect 476298 279120 476304 279132
rect 456116 279092 476304 279120
rect 456116 279080 456122 279092
rect 476298 279080 476304 279092
rect 476356 279080 476362 279132
rect 478138 279080 478144 279132
rect 478196 279120 478202 279132
rect 502702 279120 502708 279132
rect 478196 279092 502708 279120
rect 478196 279080 478202 279092
rect 502702 279080 502708 279092
rect 502760 279080 502766 279132
rect 504358 279080 504364 279132
rect 504416 279120 504422 279132
rect 518066 279120 518072 279132
rect 504416 279092 518072 279120
rect 504416 279080 504422 279092
rect 518066 279080 518072 279092
rect 518124 279080 518130 279132
rect 518158 279080 518164 279132
rect 518216 279120 518222 279132
rect 529934 279120 529940 279132
rect 518216 279092 529940 279120
rect 518216 279080 518222 279092
rect 529934 279080 529940 279092
rect 529992 279080 529998 279132
rect 87598 279012 87604 279064
rect 87656 279052 87662 279064
rect 203702 279052 203708 279064
rect 87656 279024 203708 279052
rect 87656 279012 87662 279024
rect 203702 279012 203708 279024
rect 203760 279012 203766 279064
rect 388438 279012 388444 279064
rect 388496 279052 388502 279064
rect 440510 279052 440516 279064
rect 388496 279024 440516 279052
rect 388496 279012 388502 279024
rect 440510 279012 440516 279024
rect 440568 279012 440574 279064
rect 443914 279052 443920 279064
rect 441586 279024 443920 279052
rect 86218 278944 86224 278996
rect 86276 278984 86282 278996
rect 198734 278984 198740 278996
rect 86276 278956 198740 278984
rect 86276 278944 86282 278956
rect 198734 278944 198740 278956
rect 198792 278944 198798 278996
rect 391842 278944 391848 278996
rect 391900 278984 391906 278996
rect 441586 278984 441614 279024
rect 443914 279012 443920 279024
rect 443972 279012 443978 279064
rect 460198 279012 460204 279064
rect 460256 279052 460262 279064
rect 483934 279052 483940 279064
rect 460256 279024 483940 279052
rect 460256 279012 460262 279024
rect 483934 279012 483940 279024
rect 483992 279012 483998 279064
rect 497458 279012 497464 279064
rect 497516 279052 497522 279064
rect 515490 279052 515496 279064
rect 497516 279024 515496 279052
rect 497516 279012 497522 279024
rect 515490 279012 515496 279024
rect 515548 279012 515554 279064
rect 521562 279012 521568 279064
rect 521620 279052 521626 279064
rect 527545 279055 527603 279061
rect 527545 279052 527557 279055
rect 521620 279024 527557 279052
rect 521620 279012 521626 279024
rect 527545 279021 527557 279024
rect 527591 279021 527603 279055
rect 527545 279015 527603 279021
rect 391900 278956 441614 278984
rect 391900 278944 391906 278956
rect 442258 278944 442264 278996
rect 442316 278984 442322 278996
rect 446490 278984 446496 278996
rect 442316 278956 446496 278984
rect 442316 278944 442322 278956
rect 446490 278944 446496 278956
rect 446548 278944 446554 278996
rect 468478 278944 468484 278996
rect 468536 278984 468542 278996
rect 474734 278984 474740 278996
rect 468536 278956 474740 278984
rect 468536 278944 468542 278956
rect 474734 278944 474740 278956
rect 474792 278944 474798 278996
rect 476758 278944 476764 278996
rect 476816 278984 476822 278996
rect 500126 278984 500132 278996
rect 476816 278956 500132 278984
rect 476816 278944 476822 278956
rect 500126 278944 500132 278956
rect 500184 278944 500190 278996
rect 508498 278944 508504 278996
rect 508556 278984 508562 278996
rect 521654 278984 521660 278996
rect 508556 278956 521660 278984
rect 508556 278944 508562 278956
rect 521654 278944 521660 278956
rect 521712 278944 521718 278996
rect 106918 278876 106924 278928
rect 106976 278916 106982 278928
rect 213914 278916 213920 278928
rect 106976 278888 213920 278916
rect 106976 278876 106982 278888
rect 213914 278876 213920 278888
rect 213972 278876 213978 278928
rect 409138 278876 409144 278928
rect 409196 278916 409202 278928
rect 455874 278916 455880 278928
rect 409196 278888 455880 278916
rect 409196 278876 409202 278888
rect 455874 278876 455880 278888
rect 455932 278876 455938 278928
rect 462958 278876 462964 278928
rect 463016 278916 463022 278928
rect 469585 278919 469643 278925
rect 469585 278916 469597 278919
rect 463016 278888 469597 278916
rect 463016 278876 463022 278888
rect 469585 278885 469597 278888
rect 469631 278885 469643 278919
rect 469585 278879 469643 278885
rect 475378 278876 475384 278928
rect 475436 278916 475442 278928
rect 495066 278916 495072 278928
rect 475436 278888 495072 278916
rect 475436 278876 475442 278888
rect 495066 278876 495072 278888
rect 495124 278876 495130 278928
rect 512638 278876 512644 278928
rect 512696 278916 512702 278928
rect 525794 278916 525800 278928
rect 512696 278888 525800 278916
rect 512696 278876 512702 278888
rect 525794 278876 525800 278888
rect 525852 278876 525858 278928
rect 551278 278876 551284 278928
rect 551336 278916 551342 278928
rect 558914 278916 558920 278928
rect 551336 278888 558920 278916
rect 551336 278876 551342 278888
rect 558914 278876 558920 278888
rect 558972 278876 558978 278928
rect 262306 278808 262312 278860
rect 262364 278848 262370 278860
rect 265894 278848 265900 278860
rect 262364 278820 265900 278848
rect 262364 278808 262370 278820
rect 265894 278808 265900 278820
rect 265952 278808 265958 278860
rect 405642 278808 405648 278860
rect 405700 278848 405706 278860
rect 410797 278851 410855 278857
rect 410797 278848 410809 278851
rect 405700 278820 410809 278848
rect 405700 278808 405706 278820
rect 410797 278817 410809 278820
rect 410843 278817 410855 278851
rect 410797 278811 410855 278817
rect 473998 278808 474004 278860
rect 474056 278848 474062 278860
rect 490006 278848 490012 278860
rect 474056 278820 490012 278848
rect 474056 278808 474062 278820
rect 490006 278808 490012 278820
rect 490064 278808 490070 278860
rect 556798 278808 556804 278860
rect 556856 278848 556862 278860
rect 559742 278848 559748 278860
rect 556856 278820 559748 278848
rect 556856 278808 556862 278820
rect 559742 278808 559748 278820
rect 559800 278808 559806 278860
rect 562962 278808 562968 278860
rect 563020 278848 563026 278860
rect 567470 278848 567476 278860
rect 563020 278820 567476 278848
rect 563020 278808 563026 278820
rect 567470 278808 567476 278820
rect 567528 278808 567534 278860
rect 349798 278740 349804 278792
rect 349856 278780 349862 278792
rect 354674 278780 354680 278792
rect 349856 278752 354680 278780
rect 349856 278740 349862 278752
rect 354674 278740 354680 278752
rect 354732 278740 354738 278792
rect 363598 278740 363604 278792
rect 363656 278780 363662 278792
rect 364702 278780 364708 278792
rect 363656 278752 364708 278780
rect 363656 278740 363662 278752
rect 364702 278740 364708 278752
rect 364760 278740 364766 278792
rect 383010 278740 383016 278792
rect 383068 278780 383074 278792
rect 384298 278780 384304 278792
rect 383068 278752 384304 278780
rect 383068 278740 383074 278752
rect 384298 278740 384304 278752
rect 384356 278740 384362 278792
rect 420178 278740 420184 278792
rect 420236 278780 420242 278792
rect 422662 278780 422668 278792
rect 420236 278752 422668 278780
rect 420236 278740 420242 278752
rect 422662 278740 422668 278752
rect 422720 278740 422726 278792
rect 436738 278740 436744 278792
rect 436796 278780 436802 278792
rect 441614 278780 441620 278792
rect 436796 278752 441620 278780
rect 436796 278740 436802 278752
rect 441614 278740 441620 278752
rect 441672 278740 441678 278792
rect 469858 278740 469864 278792
rect 469916 278780 469922 278792
rect 479702 278780 479708 278792
rect 469916 278752 479708 278780
rect 469916 278740 469922 278752
rect 479702 278740 479708 278752
rect 479760 278740 479766 278792
rect 555418 278740 555424 278792
rect 555476 278780 555482 278792
rect 557534 278780 557540 278792
rect 555476 278752 557540 278780
rect 555476 278740 555482 278752
rect 557534 278740 557540 278752
rect 557592 278740 557598 278792
rect 566458 278740 566464 278792
rect 566516 278780 566522 278792
rect 569126 278780 569132 278792
rect 566516 278752 569132 278780
rect 566516 278740 566522 278752
rect 569126 278740 569132 278752
rect 569184 278740 569190 278792
rect 575382 278740 575388 278792
rect 575440 278780 575446 278792
rect 576946 278780 576952 278792
rect 575440 278752 576952 278780
rect 575440 278740 575446 278752
rect 576946 278740 576952 278752
rect 577004 278740 577010 278792
rect 115198 278672 115204 278724
rect 115256 278712 115262 278724
rect 243722 278712 243728 278724
rect 115256 278684 243728 278712
rect 115256 278672 115262 278684
rect 243722 278672 243728 278684
rect 243780 278672 243786 278724
rect 278038 278672 278044 278724
rect 278096 278712 278102 278724
rect 351086 278712 351092 278724
rect 278096 278684 351092 278712
rect 278096 278672 278102 278684
rect 351086 278672 351092 278684
rect 351144 278672 351150 278724
rect 364242 278672 364248 278724
rect 364300 278712 364306 278724
rect 424226 278712 424232 278724
rect 364300 278684 424232 278712
rect 364300 278672 364306 278684
rect 424226 278672 424232 278684
rect 424284 278672 424290 278724
rect 424318 278672 424324 278724
rect 424376 278712 424382 278724
rect 465258 278712 465264 278724
rect 424376 278684 465264 278712
rect 424376 278672 424382 278684
rect 465258 278672 465264 278684
rect 465316 278672 465322 278724
rect 39298 278604 39304 278656
rect 39356 278644 39362 278656
rect 172146 278644 172152 278656
rect 39356 278616 172152 278644
rect 39356 278604 39362 278616
rect 172146 278604 172152 278616
rect 172204 278604 172210 278656
rect 291838 278604 291844 278656
rect 291896 278644 291902 278656
rect 366450 278644 366456 278656
rect 291896 278616 366456 278644
rect 291896 278604 291902 278616
rect 366450 278604 366456 278616
rect 366508 278604 366514 278656
rect 367738 278604 367744 278656
rect 367796 278644 367802 278656
rect 426894 278644 426900 278656
rect 367796 278616 426900 278644
rect 367796 278604 367802 278616
rect 426894 278604 426900 278616
rect 426952 278604 426958 278656
rect 447778 278604 447784 278656
rect 447836 278644 447842 278656
rect 481634 278644 481640 278656
rect 447836 278616 481640 278644
rect 447836 278604 447842 278616
rect 481634 278604 481640 278616
rect 481692 278604 481698 278656
rect 99282 278536 99288 278588
rect 99340 278576 99346 278588
rect 233142 278576 233148 278588
rect 99340 278548 233148 278576
rect 99340 278536 99346 278548
rect 233142 278536 233148 278548
rect 233200 278536 233206 278588
rect 289078 278536 289084 278588
rect 289136 278576 289142 278588
rect 368934 278576 368940 278588
rect 289136 278548 368940 278576
rect 289136 278536 289142 278548
rect 368934 278536 368940 278548
rect 368992 278536 368998 278588
rect 375282 278536 375288 278588
rect 375340 278576 375346 278588
rect 432046 278576 432052 278588
rect 375340 278548 432052 278576
rect 375340 278536 375346 278548
rect 432046 278536 432052 278548
rect 432104 278536 432110 278588
rect 435358 278536 435364 278588
rect 435416 278576 435422 278588
rect 475470 278576 475476 278588
rect 435416 278548 475476 278576
rect 435416 278536 435422 278548
rect 475470 278536 475476 278548
rect 475528 278536 475534 278588
rect 495894 278576 495900 278588
rect 489886 278548 495900 278576
rect 32398 278468 32404 278520
rect 32456 278508 32462 278520
rect 167914 278508 167920 278520
rect 32456 278480 167920 278508
rect 32456 278468 32462 278480
rect 167914 278468 167920 278480
rect 167972 278468 167978 278520
rect 209038 278468 209044 278520
rect 209096 278508 209102 278520
rect 293954 278508 293960 278520
rect 209096 278480 293960 278508
rect 209096 278468 209102 278480
rect 293954 278468 293960 278480
rect 294012 278468 294018 278520
rect 314010 278468 314016 278520
rect 314068 278508 314074 278520
rect 379146 278508 379152 278520
rect 314068 278480 379152 278508
rect 314068 278468 314074 278480
rect 379146 278468 379152 278480
rect 379204 278468 379210 278520
rect 382918 278468 382924 278520
rect 382976 278508 382982 278520
rect 437106 278508 437112 278520
rect 382976 278480 437112 278508
rect 382976 278468 382982 278480
rect 437106 278468 437112 278480
rect 437164 278468 437170 278520
rect 440878 278468 440884 278520
rect 440936 278508 440942 278520
rect 478046 278508 478052 278520
rect 440936 278480 478052 278508
rect 440936 278468 440942 278480
rect 478046 278468 478052 278480
rect 478104 278468 478110 278520
rect 486418 278468 486424 278520
rect 486476 278508 486482 278520
rect 489886 278508 489914 278548
rect 495894 278536 495900 278548
rect 495952 278536 495958 278588
rect 493502 278508 493508 278520
rect 486476 278480 489914 278508
rect 491772 278480 493508 278508
rect 486476 278468 486482 278480
rect 95050 278400 95056 278452
rect 95108 278440 95114 278452
rect 230934 278440 230940 278452
rect 95108 278412 230940 278440
rect 95108 278400 95114 278412
rect 230934 278400 230940 278412
rect 230992 278400 230998 278452
rect 271138 278400 271144 278452
rect 271196 278440 271202 278452
rect 355318 278440 355324 278452
rect 271196 278412 355324 278440
rect 271196 278400 271202 278412
rect 355318 278400 355324 278412
rect 355376 278400 355382 278452
rect 360102 278400 360108 278452
rect 360160 278440 360166 278452
rect 421742 278440 421748 278452
rect 360160 278412 421748 278440
rect 360160 278400 360166 278412
rect 421742 278400 421748 278412
rect 421800 278400 421806 278452
rect 425790 278400 425796 278452
rect 425848 278440 425854 278452
rect 467834 278440 467840 278452
rect 425848 278412 467840 278440
rect 425848 278400 425854 278412
rect 467834 278400 467840 278412
rect 467892 278400 467898 278452
rect 485038 278400 485044 278452
rect 485096 278440 485102 278452
rect 491772 278440 491800 278480
rect 493502 278468 493508 278480
rect 493560 278468 493566 278520
rect 485096 278412 491800 278440
rect 485096 278400 485102 278412
rect 493410 278400 493416 278452
rect 493468 278440 493474 278452
rect 503714 278440 503720 278452
rect 493468 278412 503720 278440
rect 493468 278400 493474 278412
rect 503714 278400 503720 278412
rect 503772 278400 503778 278452
rect 88978 278332 88984 278384
rect 89036 278372 89042 278384
rect 225874 278372 225880 278384
rect 89036 278344 225880 278372
rect 89036 278332 89042 278344
rect 225874 278332 225880 278344
rect 225932 278332 225938 278384
rect 258718 278332 258724 278384
rect 258776 278372 258782 278384
rect 343634 278372 343640 278384
rect 258776 278344 343640 278372
rect 258776 278332 258782 278344
rect 343634 278332 343640 278344
rect 343692 278332 343698 278384
rect 357342 278332 357348 278384
rect 357400 278372 357406 278384
rect 419534 278372 419540 278384
rect 357400 278344 419540 278372
rect 357400 278332 357406 278344
rect 419534 278332 419540 278344
rect 419592 278332 419598 278384
rect 428458 278332 428464 278384
rect 428516 278372 428522 278384
rect 470594 278372 470600 278384
rect 428516 278344 470600 278372
rect 428516 278332 428522 278344
rect 470594 278332 470600 278344
rect 470652 278332 470658 278384
rect 482278 278332 482284 278384
rect 482336 278372 482342 278384
rect 508682 278372 508688 278384
rect 482336 278344 508688 278372
rect 482336 278332 482342 278344
rect 508682 278332 508688 278344
rect 508740 278332 508746 278384
rect 25498 278264 25504 278316
rect 25556 278304 25562 278316
rect 164510 278304 164516 278316
rect 25556 278276 164516 278304
rect 25556 278264 25562 278276
rect 164510 278264 164516 278276
rect 164568 278264 164574 278316
rect 224862 278264 224868 278316
rect 224920 278304 224926 278316
rect 242802 278304 242808 278316
rect 224920 278276 242808 278304
rect 224920 278264 224926 278276
rect 242802 278264 242808 278276
rect 242860 278264 242866 278316
rect 260098 278264 260104 278316
rect 260156 278304 260162 278316
rect 348510 278304 348516 278316
rect 260156 278276 348516 278304
rect 260156 278264 260162 278276
rect 348510 278264 348516 278276
rect 348568 278264 348574 278316
rect 353938 278264 353944 278316
rect 353996 278304 354002 278316
rect 416774 278304 416780 278316
rect 353996 278276 416780 278304
rect 353996 278264 354002 278276
rect 416774 278264 416780 278276
rect 416832 278264 416838 278316
rect 417418 278264 417424 278316
rect 417476 278304 417482 278316
rect 462682 278304 462688 278316
rect 417476 278276 462688 278304
rect 417476 278264 417482 278276
rect 462682 278264 462688 278276
rect 462740 278264 462746 278316
rect 484302 278264 484308 278316
rect 484360 278304 484366 278316
rect 511258 278304 511264 278316
rect 484360 278276 511264 278304
rect 484360 278264 484366 278276
rect 511258 278264 511264 278276
rect 511316 278264 511322 278316
rect 81342 278196 81348 278248
rect 81400 278236 81406 278248
rect 220814 278236 220820 278248
rect 81400 278208 220820 278236
rect 81400 278196 81406 278208
rect 220814 278196 220820 278208
rect 220872 278196 220878 278248
rect 242158 278196 242164 278248
rect 242216 278236 242222 278248
rect 332594 278236 332600 278248
rect 242216 278208 332600 278236
rect 242216 278196 242222 278208
rect 332594 278196 332600 278208
rect 332652 278196 332658 278248
rect 342070 278196 342076 278248
rect 342128 278236 342134 278248
rect 409046 278236 409052 278248
rect 342128 278208 409052 278236
rect 342128 278196 342134 278208
rect 409046 278196 409052 278208
rect 409104 278196 409110 278248
rect 410518 278196 410524 278248
rect 410576 278236 410582 278248
rect 457530 278236 457536 278248
rect 410576 278208 457536 278236
rect 410576 278196 410582 278208
rect 457530 278196 457536 278208
rect 457588 278196 457594 278248
rect 471238 278196 471244 278248
rect 471296 278236 471302 278248
rect 501046 278236 501052 278248
rect 471296 278208 501052 278236
rect 471296 278196 471302 278208
rect 501046 278196 501052 278208
rect 501104 278196 501110 278248
rect 22738 278128 22744 278180
rect 22796 278168 22802 278180
rect 163682 278168 163688 278180
rect 22796 278140 163688 278168
rect 22796 278128 22802 278140
rect 163682 278128 163688 278140
rect 163740 278128 163746 278180
rect 240778 278128 240784 278180
rect 240836 278168 240842 278180
rect 333146 278168 333152 278180
rect 240836 278140 333152 278168
rect 240836 278128 240842 278140
rect 333146 278128 333152 278140
rect 333204 278128 333210 278180
rect 339402 278128 339408 278180
rect 339460 278168 339466 278180
rect 406470 278168 406476 278180
rect 339460 278140 406476 278168
rect 339460 278128 339466 278140
rect 406470 278128 406476 278140
rect 406528 278128 406534 278180
rect 407022 278128 407028 278180
rect 407080 278168 407086 278180
rect 455046 278168 455052 278180
rect 407080 278140 455052 278168
rect 407080 278128 407086 278140
rect 455046 278128 455052 278140
rect 455104 278128 455110 278180
rect 466270 278128 466276 278180
rect 466328 278168 466334 278180
rect 498470 278168 498476 278180
rect 466328 278140 498476 278168
rect 466328 278128 466334 278140
rect 498470 278128 498476 278140
rect 498528 278128 498534 278180
rect 48222 278060 48228 278112
rect 48280 278100 48286 278112
rect 196894 278100 196900 278112
rect 48280 278072 196900 278100
rect 48280 278060 48286 278072
rect 196894 278060 196900 278072
rect 196952 278060 196958 278112
rect 233142 278060 233148 278112
rect 233200 278100 233206 278112
rect 329834 278100 329840 278112
rect 233200 278072 329840 278100
rect 233200 278060 233206 278072
rect 329834 278060 329840 278072
rect 329892 278060 329898 278112
rect 331858 278060 331864 278112
rect 331916 278100 331922 278112
rect 399662 278100 399668 278112
rect 331916 278072 399668 278100
rect 331916 278060 331922 278072
rect 399662 278060 399668 278072
rect 399720 278060 399726 278112
rect 400858 278060 400864 278112
rect 400916 278100 400922 278112
rect 449894 278100 449900 278112
rect 400916 278072 449900 278100
rect 400916 278060 400922 278072
rect 449894 278060 449900 278072
rect 449952 278060 449958 278112
rect 450538 278060 450544 278112
rect 450596 278100 450602 278112
rect 485774 278100 485780 278112
rect 450596 278072 485780 278100
rect 450596 278060 450602 278072
rect 485774 278060 485780 278072
rect 485832 278060 485838 278112
rect 489178 278060 489184 278112
rect 489236 278100 489242 278112
rect 513742 278100 513748 278112
rect 489236 278072 513748 278100
rect 489236 278060 489242 278072
rect 513742 278060 513748 278072
rect 513800 278060 513806 278112
rect 14458 277992 14464 278044
rect 14516 278032 14522 278044
rect 162854 278032 162860 278044
rect 14516 278004 162860 278032
rect 14516 277992 14522 278004
rect 162854 277992 162860 278004
rect 162912 277992 162918 278044
rect 227622 277992 227628 278044
rect 227680 278032 227686 278044
rect 325878 278032 325884 278044
rect 227680 278004 325884 278032
rect 227680 277992 227686 278004
rect 325878 277992 325884 278004
rect 325936 277992 325942 278044
rect 332502 277992 332508 278044
rect 332560 278032 332566 278044
rect 401594 278032 401600 278044
rect 332560 278004 401600 278032
rect 332560 277992 332566 278004
rect 401594 277992 401600 278004
rect 401652 277992 401658 278044
rect 403618 277992 403624 278044
rect 403676 278032 403682 278044
rect 452654 278032 452660 278044
rect 403676 278004 452660 278032
rect 403676 277992 403682 278004
rect 452654 277992 452660 278004
rect 452712 277992 452718 278044
rect 453298 277992 453304 278044
rect 453356 278032 453362 278044
rect 488534 278032 488540 278044
rect 453356 278004 488540 278032
rect 453356 277992 453362 278004
rect 488534 277992 488540 278004
rect 488592 277992 488598 278044
rect 491202 277992 491208 278044
rect 491260 278032 491266 278044
rect 516318 278032 516324 278044
rect 491260 278004 516324 278032
rect 491260 277992 491266 278004
rect 516318 277992 516324 278004
rect 516376 277992 516382 278044
rect 135162 277924 135168 277976
rect 135220 277964 135226 277976
rect 259086 277964 259092 277976
rect 135220 277936 259092 277964
rect 135220 277924 135226 277936
rect 259086 277924 259092 277936
rect 259144 277924 259150 277976
rect 316678 277924 316684 277976
rect 316736 277964 316742 277976
rect 374086 277964 374092 277976
rect 316736 277936 374092 277964
rect 316736 277924 316742 277936
rect 374086 277924 374092 277936
rect 374144 277924 374150 277976
rect 392578 277924 392584 277976
rect 392636 277964 392642 277976
rect 444742 277964 444748 277976
rect 392636 277936 444748 277964
rect 392636 277924 392642 277936
rect 444742 277924 444748 277936
rect 444800 277924 444806 277976
rect 446398 277924 446404 277976
rect 446456 277964 446462 277976
rect 480530 277964 480536 277976
rect 446456 277936 480536 277964
rect 446456 277924 446462 277936
rect 480530 277924 480536 277936
rect 480588 277924 480594 277976
rect 151722 277856 151728 277908
rect 151780 277896 151786 277908
rect 270954 277896 270960 277908
rect 151780 277868 270960 277896
rect 151780 277856 151786 277868
rect 270954 277856 270960 277868
rect 271012 277856 271018 277908
rect 335998 277856 336004 277908
rect 336056 277896 336062 277908
rect 386874 277896 386880 277908
rect 336056 277868 386880 277896
rect 336056 277856 336062 277868
rect 386874 277856 386880 277868
rect 386932 277856 386938 277908
rect 389910 277856 389916 277908
rect 389968 277896 389974 277908
rect 442350 277896 442356 277908
rect 389968 277868 442356 277896
rect 389968 277856 389974 277868
rect 442350 277856 442356 277868
rect 442408 277856 442414 277908
rect 144822 277788 144828 277840
rect 144880 277828 144886 277840
rect 262306 277828 262312 277840
rect 144880 277800 262312 277828
rect 144880 277788 144886 277800
rect 262306 277788 262312 277800
rect 262364 277788 262370 277840
rect 396718 277788 396724 277840
rect 396776 277828 396782 277840
rect 447318 277828 447324 277840
rect 396776 277800 447324 277828
rect 396776 277788 396782 277800
rect 447318 277788 447324 277800
rect 447376 277788 447382 277840
rect 246298 277720 246304 277772
rect 246356 277760 246362 277772
rect 311894 277760 311900 277772
rect 246356 277732 311900 277760
rect 246356 277720 246362 277732
rect 311894 277720 311900 277732
rect 311952 277720 311958 277772
rect 413922 277720 413928 277772
rect 413980 277760 413986 277772
rect 460106 277760 460112 277772
rect 413980 277732 460112 277760
rect 413980 277720 413986 277732
rect 460106 277720 460112 277732
rect 460164 277720 460170 277772
rect 231118 277652 231124 277704
rect 231176 277692 231182 277704
rect 296714 277692 296720 277704
rect 231176 277664 296720 277692
rect 231176 277652 231182 277664
rect 296714 277652 296720 277664
rect 296772 277652 296778 277704
rect 250438 277584 250444 277636
rect 250496 277624 250502 277636
rect 314654 277624 314660 277636
rect 250496 277596 314660 277624
rect 250496 277584 250502 277596
rect 314654 277584 314660 277596
rect 314712 277584 314718 277636
rect 238018 277516 238024 277568
rect 238076 277556 238082 277568
rect 301682 277556 301688 277568
rect 238076 277528 301688 277556
rect 238076 277516 238082 277528
rect 301682 277516 301688 277528
rect 301740 277516 301746 277568
rect 262858 277448 262864 277500
rect 262916 277488 262922 277500
rect 319530 277488 319536 277500
rect 262916 277460 319536 277488
rect 262916 277448 262922 277460
rect 319530 277448 319536 277460
rect 319588 277448 319594 277500
rect 253198 277380 253204 277432
rect 253256 277420 253262 277432
rect 299106 277420 299112 277432
rect 253256 277392 299112 277420
rect 253256 277380 253262 277392
rect 299106 277380 299112 277392
rect 299164 277380 299170 277432
rect 137922 277312 137928 277364
rect 137980 277352 137986 277364
rect 255406 277352 255412 277364
rect 137980 277324 255412 277352
rect 137980 277312 137986 277324
rect 255406 277312 255412 277324
rect 255464 277312 255470 277364
rect 153102 277244 153108 277296
rect 153160 277284 153166 277296
rect 271782 277284 271788 277296
rect 153160 277256 271788 277284
rect 153160 277244 153166 277256
rect 271782 277244 271788 277256
rect 271840 277244 271846 277296
rect 273898 277244 273904 277296
rect 273956 277284 273962 277296
rect 340966 277284 340972 277296
rect 273956 277256 340972 277284
rect 273956 277244 273962 277256
rect 340966 277244 340972 277256
rect 341024 277244 341030 277296
rect 155862 277176 155868 277228
rect 155920 277216 155926 277228
rect 274542 277216 274548 277228
rect 155920 277188 274548 277216
rect 155920 277176 155926 277188
rect 274542 277176 274548 277188
rect 274600 277176 274606 277228
rect 112438 277108 112444 277160
rect 112496 277148 112502 277160
rect 240226 277148 240232 277160
rect 112496 277120 240232 277148
rect 112496 277108 112502 277120
rect 240226 277108 240232 277120
rect 240284 277108 240290 277160
rect 266998 277108 267004 277160
rect 267056 277148 267062 277160
rect 338206 277148 338212 277160
rect 267056 277120 338212 277148
rect 267056 277108 267062 277120
rect 338206 277108 338212 277120
rect 338264 277108 338270 277160
rect 347038 277108 347044 277160
rect 347096 277148 347102 277160
rect 401778 277148 401784 277160
rect 347096 277120 401784 277148
rect 347096 277108 347102 277120
rect 401778 277108 401784 277120
rect 401836 277108 401842 277160
rect 105538 277040 105544 277092
rect 105596 277080 105602 277092
rect 236086 277080 236092 277092
rect 105596 277052 236092 277080
rect 105596 277040 105602 277052
rect 236086 277040 236092 277052
rect 236144 277040 236150 277092
rect 280798 277040 280804 277092
rect 280856 277080 280862 277092
rect 356146 277080 356152 277092
rect 280856 277052 356152 277080
rect 280856 277040 280862 277052
rect 356146 277040 356152 277052
rect 356204 277040 356210 277092
rect 54478 276972 54484 277024
rect 54536 277012 54542 277024
rect 185026 277012 185032 277024
rect 54536 276984 185032 277012
rect 54536 276972 54542 276984
rect 185026 276972 185032 276984
rect 185084 276972 185090 277024
rect 284938 276972 284944 277024
rect 284996 277012 285002 277024
rect 361574 277012 361580 277024
rect 284996 276984 361580 277012
rect 284996 276972 285002 276984
rect 361574 276972 361580 276984
rect 361632 276972 361638 277024
rect 106182 276904 106188 276956
rect 106240 276944 106246 276956
rect 238662 276944 238668 276956
rect 106240 276916 238668 276944
rect 106240 276904 106246 276916
rect 238662 276904 238668 276916
rect 238720 276904 238726 276956
rect 286318 276904 286324 276956
rect 286376 276944 286382 276956
rect 363046 276944 363052 276956
rect 286376 276916 363052 276944
rect 286376 276904 286382 276916
rect 363046 276904 363052 276916
rect 363104 276904 363110 276956
rect 58618 276836 58624 276888
rect 58676 276876 58682 276888
rect 191926 276876 191932 276888
rect 58676 276848 191932 276876
rect 58676 276836 58682 276848
rect 191926 276836 191932 276848
rect 191984 276836 191990 276888
rect 220722 276836 220728 276888
rect 220780 276876 220786 276888
rect 317506 276876 317512 276888
rect 220780 276848 317512 276876
rect 220780 276836 220786 276848
rect 317506 276836 317512 276848
rect 317564 276836 317570 276888
rect 324958 276836 324964 276888
rect 325016 276876 325022 276888
rect 394786 276876 394792 276888
rect 325016 276848 394792 276876
rect 325016 276836 325022 276848
rect 394786 276836 394792 276848
rect 394844 276836 394850 276888
rect 93118 276768 93124 276820
rect 93176 276808 93182 276820
rect 227990 276808 227996 276820
rect 93176 276780 227996 276808
rect 93176 276768 93182 276780
rect 227990 276768 227996 276780
rect 228048 276768 228054 276820
rect 282178 276768 282184 276820
rect 282236 276808 282242 276820
rect 358906 276808 358912 276820
rect 282236 276780 358912 276808
rect 282236 276768 282242 276780
rect 358906 276768 358912 276780
rect 358964 276768 358970 276820
rect 360838 276768 360844 276820
rect 360896 276808 360902 276820
rect 404354 276808 404360 276820
rect 360896 276780 404360 276808
rect 360896 276768 360902 276780
rect 404354 276768 404360 276780
rect 404412 276768 404418 276820
rect 40678 276700 40684 276752
rect 40736 276740 40742 276752
rect 178126 276740 178132 276752
rect 40736 276712 178132 276740
rect 40736 276700 40742 276712
rect 178126 276700 178132 276712
rect 178184 276700 178190 276752
rect 227530 276700 227536 276752
rect 227588 276740 227594 276752
rect 325602 276740 325608 276752
rect 227588 276712 325608 276740
rect 227588 276700 227594 276712
rect 325602 276700 325608 276712
rect 325660 276700 325666 276752
rect 340138 276700 340144 276752
rect 340196 276740 340202 276752
rect 396166 276740 396172 276752
rect 340196 276712 396172 276740
rect 340196 276700 340202 276712
rect 396166 276700 396172 276712
rect 396224 276700 396230 276752
rect 33778 276632 33784 276684
rect 33836 276672 33842 276684
rect 175274 276672 175280 276684
rect 33836 276644 175280 276672
rect 33836 276632 33842 276644
rect 175274 276632 175280 276644
rect 175332 276632 175338 276684
rect 215938 276632 215944 276684
rect 215996 276672 216002 276684
rect 316126 276672 316132 276684
rect 215996 276644 316132 276672
rect 215996 276632 216002 276644
rect 316126 276632 316132 276644
rect 316184 276632 316190 276684
rect 318058 276632 318064 276684
rect 318116 276672 318122 276684
rect 389174 276672 389180 276684
rect 318116 276644 389180 276672
rect 318116 276632 318122 276644
rect 389174 276632 389180 276644
rect 389232 276632 389238 276684
rect 431862 276632 431868 276684
rect 431920 276672 431926 276684
rect 472066 276672 472072 276684
rect 431920 276644 472072 276672
rect 431920 276632 431926 276644
rect 472066 276632 472072 276644
rect 472124 276632 472130 276684
rect 160002 276564 160008 276616
rect 160060 276604 160066 276616
rect 276106 276604 276112 276616
rect 160060 276576 276112 276604
rect 160060 276564 160066 276576
rect 276106 276564 276112 276576
rect 276164 276564 276170 276616
rect 117222 276496 117228 276548
rect 117280 276536 117286 276548
rect 226978 276536 226984 276548
rect 117280 276508 226984 276536
rect 117280 276496 117286 276508
rect 226978 276496 226984 276508
rect 227036 276496 227042 276548
rect 51718 275408 51724 275460
rect 51776 275448 51782 275460
rect 182174 275448 182180 275460
rect 51776 275420 182180 275448
rect 51776 275408 51782 275420
rect 182174 275408 182180 275420
rect 182232 275408 182238 275460
rect 57238 275340 57244 275392
rect 57296 275380 57302 275392
rect 187786 275380 187792 275392
rect 57296 275352 187792 275380
rect 57296 275340 57302 275352
rect 187786 275340 187792 275352
rect 187844 275340 187850 275392
rect 61378 275272 61384 275324
rect 61436 275312 61442 275324
rect 194778 275312 194784 275324
rect 61436 275284 194784 275312
rect 61436 275272 61442 275284
rect 194778 275272 194784 275284
rect 194836 275272 194842 275324
rect 124122 271124 124128 271176
rect 124180 271164 124186 271176
rect 208486 271164 208492 271176
rect 124180 271136 208492 271164
rect 124180 271124 124186 271136
rect 208486 271124 208492 271136
rect 208544 271124 208550 271176
rect 161382 265616 161388 265668
rect 161440 265656 161446 265668
rect 252002 265656 252008 265668
rect 161440 265628 252008 265656
rect 161440 265616 161446 265628
rect 252002 265616 252008 265628
rect 252060 265616 252066 265668
rect 245010 259360 245016 259412
rect 245068 259400 245074 259412
rect 580166 259400 580172 259412
rect 245068 259372 580172 259400
rect 245068 259360 245074 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 3418 255212 3424 255264
rect 3476 255252 3482 255264
rect 68278 255252 68284 255264
rect 3476 255224 68284 255252
rect 3476 255212 3482 255224
rect 68278 255212 68284 255224
rect 68336 255212 68342 255264
rect 119982 254532 119988 254584
rect 120040 254572 120046 254584
rect 222838 254572 222844 254584
rect 120040 254544 222844 254572
rect 120040 254532 120046 254544
rect 222838 254532 222844 254544
rect 222896 254532 222902 254584
rect 582926 245596 582932 245608
rect 582887 245568 582932 245596
rect 582926 245556 582932 245568
rect 582984 245556 582990 245608
rect 133782 243516 133788 243568
rect 133840 243556 133846 243568
rect 258074 243556 258080 243568
rect 133840 243528 258080 243556
rect 133840 243516 133846 243528
rect 258074 243516 258080 243528
rect 258132 243516 258138 243568
rect 258810 243516 258816 243568
rect 258868 243556 258874 243568
rect 329834 243556 329840 243568
rect 258868 243528 329840 243556
rect 258868 243516 258874 243528
rect 329834 243516 329840 243528
rect 329892 243516 329898 243568
rect 3418 241408 3424 241460
rect 3476 241448 3482 241460
rect 53190 241448 53196 241460
rect 3476 241420 53196 241448
rect 3476 241408 3482 241420
rect 53190 241408 53196 241420
rect 53248 241408 53254 241460
rect 147582 238008 147588 238060
rect 147640 238048 147646 238060
rect 268010 238048 268016 238060
rect 147640 238020 268016 238048
rect 147640 238008 147646 238020
rect 268010 238008 268016 238020
rect 268068 238008 268074 238060
rect 233970 219376 233976 219428
rect 234028 219416 234034 219428
rect 579982 219416 579988 219428
rect 234028 219388 579988 219416
rect 234028 219376 234034 219388
rect 579982 219376 579988 219388
rect 580040 219376 580046 219428
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 65518 189020 65524 189032
rect 3476 188992 65524 189020
rect 3476 188980 3482 188992
rect 65518 188980 65524 188992
rect 65576 188980 65582 189032
rect 231210 179324 231216 179376
rect 231268 179364 231274 179376
rect 580166 179364 580172 179376
rect 231268 179336 580172 179364
rect 231268 179324 231274 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 148318 164200 148324 164212
rect 3292 164172 148324 164200
rect 3292 164160 3298 164172
rect 148318 164160 148324 164172
rect 148376 164160 148382 164212
rect 233970 163548 233976 163600
rect 234028 163588 234034 163600
rect 316034 163588 316040 163600
rect 234028 163560 316040 163588
rect 234028 163548 234034 163560
rect 316034 163548 316040 163560
rect 316092 163548 316098 163600
rect 148962 163480 148968 163532
rect 149020 163520 149026 163532
rect 269206 163520 269212 163532
rect 149020 163492 269212 163520
rect 149020 163480 149026 163492
rect 269206 163480 269212 163492
rect 269264 163480 269270 163532
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 71038 150396 71044 150408
rect 3476 150368 71044 150396
rect 3476 150356 3482 150368
rect 71038 150356 71044 150368
rect 71096 150356 71102 150408
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 21358 137952 21364 137964
rect 3292 137924 21364 137952
rect 3292 137912 3298 137924
rect 21358 137912 21364 137924
rect 21416 137912 21422 137964
rect 582466 126052 582472 126064
rect 582427 126024 582472 126052
rect 582466 126012 582472 126024
rect 582524 126012 582530 126064
rect 162394 113092 162400 113144
rect 162452 113132 162458 113144
rect 580166 113132 580172 113144
rect 162452 113104 580172 113132
rect 162452 113092 162458 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 141418 111772 141424 111784
rect 3476 111744 141424 111772
rect 3476 111732 3482 111744
rect 141418 111732 141424 111744
rect 141476 111732 141482 111784
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 53098 97968 53104 97980
rect 3476 97940 53104 97968
rect 3476 97928 3482 97940
rect 53098 97928 53104 97940
rect 53156 97928 53162 97980
rect 350442 93100 350448 93152
rect 350500 93140 350506 93152
rect 414106 93140 414112 93152
rect 350500 93112 414112 93140
rect 350500 93100 350506 93112
rect 414106 93100 414112 93112
rect 414164 93100 414170 93152
rect 472710 91740 472716 91792
rect 472768 91780 472774 91792
rect 490006 91780 490012 91792
rect 472768 91752 490012 91780
rect 472768 91740 472774 91752
rect 490006 91740 490012 91752
rect 490064 91740 490070 91792
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 582837 85527 582895 85533
rect 582837 85524 582849 85527
rect 3200 85496 582849 85524
rect 3200 85484 3206 85496
rect 582837 85493 582849 85496
rect 582883 85493 582895 85527
rect 582837 85487 582895 85493
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 582745 71723 582803 71729
rect 582745 71720 582757 71723
rect 3476 71692 582757 71720
rect 3476 71680 3482 71692
rect 582745 71689 582757 71692
rect 582791 71689 582803 71723
rect 582745 71683 582803 71689
rect 142062 71000 142068 71052
rect 142120 71040 142126 71052
rect 263778 71040 263784 71052
rect 142120 71012 263784 71040
rect 142120 71000 142126 71012
rect 263778 71000 263784 71012
rect 263836 71000 263842 71052
rect 162486 60664 162492 60716
rect 162544 60704 162550 60716
rect 579890 60704 579896 60716
rect 162544 60676 579896 60704
rect 162544 60664 162550 60676
rect 579890 60664 579896 60676
rect 579948 60664 579954 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 582653 59347 582711 59353
rect 582653 59344 582665 59347
rect 3108 59316 582665 59344
rect 3108 59304 3114 59316
rect 582653 59313 582665 59316
rect 582699 59313 582711 59347
rect 582653 59307 582711 59313
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 582561 45543 582619 45549
rect 582561 45540 582573 45543
rect 3476 45512 582573 45540
rect 3476 45500 3482 45512
rect 582561 45509 582573 45512
rect 582607 45509 582619 45543
rect 582561 45503 582619 45509
rect 255958 36524 255964 36576
rect 256016 36564 256022 36576
rect 303798 36564 303804 36576
rect 256016 36536 303804 36564
rect 256016 36524 256022 36536
rect 303798 36524 303804 36536
rect 303856 36524 303862 36576
rect 162578 33056 162584 33108
rect 162636 33096 162642 33108
rect 580166 33096 580172 33108
rect 162636 33068 580172 33096
rect 162636 33056 162642 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 162670 20612 162676 20664
rect 162728 20652 162734 20664
rect 580166 20652 580172 20664
rect 162728 20624 580172 20652
rect 162728 20612 162734 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 129642 17212 129648 17264
rect 129700 17252 129706 17264
rect 255314 17252 255320 17264
rect 129700 17224 255320 17252
rect 129700 17212 129706 17224
rect 255314 17212 255320 17224
rect 255372 17212 255378 17264
rect 126882 13064 126888 13116
rect 126940 13104 126946 13116
rect 252738 13104 252744 13116
rect 126940 13076 252744 13104
rect 126940 13064 126946 13076
rect 252738 13064 252744 13076
rect 252796 13064 252802 13116
rect 245010 12112 245016 12164
rect 245068 12152 245074 12164
rect 306374 12152 306380 12164
rect 245068 12124 306380 12152
rect 245068 12112 245074 12124
rect 306374 12112 306380 12124
rect 306432 12112 306438 12164
rect 228634 12044 228640 12096
rect 228692 12084 228698 12096
rect 324314 12084 324320 12096
rect 228692 12056 324320 12084
rect 228692 12044 228698 12056
rect 324314 12044 324320 12056
rect 324372 12044 324378 12096
rect 230934 11976 230940 12028
rect 230992 12016 230998 12028
rect 327166 12016 327172 12028
rect 230992 11988 327172 12016
rect 230992 11976 230998 11988
rect 327166 11976 327172 11988
rect 327224 11976 327230 12028
rect 224218 11908 224224 11960
rect 224276 11948 224282 11960
rect 321738 11948 321744 11960
rect 224276 11920 321744 11948
rect 224276 11908 224282 11920
rect 321738 11908 321744 11920
rect 321796 11908 321802 11960
rect 223482 11840 223488 11892
rect 223540 11880 223546 11892
rect 323026 11880 323032 11892
rect 223540 11852 323032 11880
rect 223540 11840 223546 11852
rect 323026 11840 323032 11852
rect 323084 11840 323090 11892
rect 342070 11840 342076 11892
rect 342128 11840 342134 11892
rect 158622 11772 158628 11824
rect 158680 11812 158686 11824
rect 276014 11812 276020 11824
rect 158680 11784 276020 11812
rect 158680 11772 158686 11784
rect 276014 11772 276020 11784
rect 276072 11772 276078 11824
rect 144730 11704 144736 11756
rect 144788 11744 144794 11756
rect 266354 11744 266360 11756
rect 144788 11716 266360 11744
rect 144788 11704 144794 11716
rect 266354 11704 266360 11716
rect 266412 11704 266418 11756
rect 342088 11676 342116 11840
rect 342162 11676 342168 11688
rect 342088 11648 342168 11676
rect 342162 11636 342168 11648
rect 342220 11636 342226 11688
rect 169662 10956 169668 11008
rect 169720 10996 169726 11008
rect 244918 10996 244924 11008
rect 169720 10968 244924 10996
rect 169720 10956 169726 10968
rect 244918 10956 244924 10968
rect 244976 10956 244982 11008
rect 165522 10888 165528 10940
rect 165580 10928 165586 10940
rect 251910 10928 251916 10940
rect 165580 10900 251916 10928
rect 165580 10888 165586 10900
rect 251910 10888 251916 10900
rect 251968 10888 251974 10940
rect 179046 10820 179052 10872
rect 179104 10860 179110 10872
rect 291194 10860 291200 10872
rect 179104 10832 291200 10860
rect 179104 10820 179110 10832
rect 291194 10820 291200 10832
rect 291252 10820 291258 10872
rect 176562 10752 176568 10804
rect 176620 10792 176626 10804
rect 288526 10792 288532 10804
rect 176620 10764 288532 10792
rect 176620 10752 176626 10764
rect 288526 10752 288532 10764
rect 288584 10752 288590 10804
rect 136450 10684 136456 10736
rect 136508 10724 136514 10736
rect 249058 10724 249064 10736
rect 136508 10696 249064 10724
rect 136508 10684 136514 10696
rect 249058 10684 249064 10696
rect 249116 10684 249122 10736
rect 154206 10616 154212 10668
rect 154264 10656 154270 10668
rect 273254 10656 273260 10668
rect 154264 10628 273260 10656
rect 154264 10616 154270 10628
rect 273254 10616 273260 10628
rect 273312 10616 273318 10668
rect 140682 10548 140688 10600
rect 140740 10588 140746 10600
rect 263594 10588 263600 10600
rect 140740 10560 263600 10588
rect 140740 10548 140746 10560
rect 263594 10548 263600 10560
rect 263652 10548 263658 10600
rect 128170 10480 128176 10532
rect 128228 10520 128234 10532
rect 251818 10520 251824 10532
rect 128228 10492 251824 10520
rect 128228 10480 128234 10492
rect 251818 10480 251824 10492
rect 251876 10480 251882 10532
rect 252002 10480 252008 10532
rect 252060 10520 252066 10532
rect 309226 10520 309232 10532
rect 252060 10492 309232 10520
rect 252060 10480 252066 10492
rect 309226 10480 309232 10492
rect 309284 10480 309290 10532
rect 85482 10412 85488 10464
rect 85540 10452 85546 10464
rect 223574 10452 223580 10464
rect 85540 10424 223580 10452
rect 85540 10412 85546 10424
rect 223574 10412 223580 10424
rect 223632 10412 223638 10464
rect 268378 10412 268384 10464
rect 268436 10452 268442 10464
rect 353294 10452 353300 10464
rect 268436 10424 353300 10452
rect 268436 10412 268442 10424
rect 353294 10412 353300 10424
rect 353352 10412 353358 10464
rect 162762 10344 162768 10396
rect 162820 10384 162826 10396
rect 580258 10384 580264 10396
rect 162820 10356 580264 10384
rect 162820 10344 162826 10356
rect 580258 10344 580264 10356
rect 580316 10344 580322 10396
rect 3418 10276 3424 10328
rect 3476 10316 3482 10328
rect 582377 10319 582435 10325
rect 582377 10316 582389 10319
rect 3476 10288 582389 10316
rect 3476 10276 3482 10288
rect 582377 10285 582389 10288
rect 582423 10285 582435 10319
rect 582377 10279 582435 10285
rect 149514 9596 149520 9648
rect 149572 9636 149578 9648
rect 269114 9636 269120 9648
rect 149572 9608 269120 9636
rect 149572 9596 149578 9608
rect 269114 9596 269120 9608
rect 269172 9596 269178 9648
rect 153010 9528 153016 9580
rect 153068 9568 153074 9580
rect 271966 9568 271972 9580
rect 153068 9540 271972 9568
rect 153068 9528 153074 9540
rect 271966 9528 271972 9540
rect 272024 9528 272030 9580
rect 145926 9460 145932 9512
rect 145984 9500 145990 9512
rect 267734 9500 267740 9512
rect 145984 9472 267740 9500
rect 145984 9460 145990 9472
rect 267734 9460 267740 9472
rect 267792 9460 267798 9512
rect 142430 9392 142436 9444
rect 142488 9432 142494 9444
rect 265066 9432 265072 9444
rect 142488 9404 265072 9432
rect 142488 9392 142494 9404
rect 265066 9392 265072 9404
rect 265124 9392 265130 9444
rect 138842 9324 138848 9376
rect 138900 9364 138906 9376
rect 262214 9364 262220 9376
rect 138900 9336 262220 9364
rect 138900 9324 138906 9336
rect 262214 9324 262220 9336
rect 262272 9324 262278 9376
rect 122282 9256 122288 9308
rect 122340 9296 122346 9308
rect 249886 9296 249892 9308
rect 122340 9268 249892 9296
rect 122340 9256 122346 9268
rect 249886 9256 249892 9268
rect 249944 9256 249950 9308
rect 118786 9188 118792 9240
rect 118844 9228 118850 9240
rect 247126 9228 247132 9240
rect 118844 9200 247132 9228
rect 118844 9188 118850 9200
rect 247126 9188 247132 9200
rect 247184 9188 247190 9240
rect 267826 9188 267832 9240
rect 267884 9228 267890 9240
rect 335354 9228 335360 9240
rect 267884 9200 335360 9228
rect 267884 9188 267890 9200
rect 335354 9188 335360 9200
rect 335412 9188 335418 9240
rect 115290 9120 115296 9172
rect 115348 9160 115354 9172
rect 245746 9160 245752 9172
rect 115348 9132 245752 9160
rect 115348 9120 115354 9132
rect 245746 9120 245752 9132
rect 245804 9120 245810 9172
rect 269114 9120 269120 9172
rect 269172 9160 269178 9172
rect 345106 9160 345112 9172
rect 269172 9132 345112 9160
rect 269172 9120 269178 9132
rect 345106 9120 345112 9132
rect 345164 9120 345170 9172
rect 108114 9052 108120 9104
rect 108172 9092 108178 9104
rect 240134 9092 240140 9104
rect 108172 9064 240140 9092
rect 108172 9052 108178 9064
rect 240134 9052 240140 9064
rect 240192 9052 240198 9104
rect 258074 9052 258080 9104
rect 258132 9092 258138 9104
rect 342254 9092 342260 9104
rect 258132 9064 342260 9092
rect 258132 9052 258138 9064
rect 342254 9052 342260 9064
rect 342312 9052 342318 9104
rect 111610 8984 111616 9036
rect 111668 9024 111674 9036
rect 242894 9024 242900 9036
rect 111668 8996 242900 9024
rect 111668 8984 111674 8996
rect 242894 8984 242900 8996
rect 242952 8984 242958 9036
rect 264146 8984 264152 9036
rect 264204 9024 264210 9036
rect 352006 9024 352012 9036
rect 264204 8996 352012 9024
rect 264204 8984 264210 8996
rect 352006 8984 352012 8996
rect 352064 8984 352070 9036
rect 104526 8916 104532 8968
rect 104584 8956 104590 8968
rect 237374 8956 237380 8968
rect 104584 8928 237380 8956
rect 104584 8916 104590 8928
rect 237374 8916 237380 8928
rect 237432 8916 237438 8968
rect 240134 8916 240140 8968
rect 240192 8956 240198 8968
rect 334066 8956 334072 8968
rect 240192 8928 334072 8956
rect 240192 8916 240198 8928
rect 334066 8916 334072 8928
rect 334124 8916 334130 8968
rect 156598 8848 156604 8900
rect 156656 8888 156662 8900
rect 274910 8888 274916 8900
rect 156656 8860 274916 8888
rect 156656 8848 156662 8860
rect 274910 8848 274916 8860
rect 274968 8848 274974 8900
rect 160094 8780 160100 8832
rect 160152 8820 160158 8832
rect 277394 8820 277400 8832
rect 160152 8792 277400 8820
rect 160152 8780 160158 8792
rect 277394 8780 277400 8792
rect 277452 8780 277458 8832
rect 171962 8712 171968 8764
rect 172020 8752 172026 8764
rect 233878 8752 233884 8764
rect 172020 8724 233884 8752
rect 172020 8712 172026 8724
rect 233878 8712 233884 8724
rect 233936 8712 233942 8764
rect 233970 8712 233976 8764
rect 234028 8752 234034 8764
rect 327074 8752 327080 8764
rect 234028 8724 327080 8752
rect 234028 8712 234034 8724
rect 327074 8712 327080 8724
rect 327132 8712 327138 8764
rect 237374 8644 237380 8696
rect 237432 8684 237438 8696
rect 320174 8684 320180 8696
rect 237432 8656 320180 8684
rect 237432 8644 237438 8656
rect 320174 8644 320180 8656
rect 320232 8644 320238 8696
rect 177850 8236 177856 8288
rect 177908 8276 177914 8288
rect 289906 8276 289912 8288
rect 177908 8248 289912 8276
rect 177908 8236 177914 8248
rect 289906 8236 289912 8248
rect 289964 8236 289970 8288
rect 167178 8168 167184 8220
rect 167236 8208 167242 8220
rect 283006 8208 283012 8220
rect 167236 8180 283012 8208
rect 167236 8168 167242 8180
rect 283006 8168 283012 8180
rect 283064 8168 283070 8220
rect 170766 8100 170772 8152
rect 170824 8140 170830 8152
rect 285766 8140 285772 8152
rect 170824 8112 285772 8140
rect 170824 8100 170830 8112
rect 285766 8100 285772 8112
rect 285824 8100 285830 8152
rect 163682 8032 163688 8084
rect 163740 8072 163746 8084
rect 280154 8072 280160 8084
rect 163740 8044 280160 8072
rect 163740 8032 163746 8044
rect 280154 8032 280160 8044
rect 280212 8032 280218 8084
rect 135254 7964 135260 8016
rect 135312 8004 135318 8016
rect 259546 8004 259552 8016
rect 135312 7976 259552 8004
rect 135312 7964 135318 7976
rect 259546 7964 259552 7976
rect 259604 7964 259610 8016
rect 131758 7896 131764 7948
rect 131816 7936 131822 7948
rect 256970 7936 256976 7948
rect 131816 7908 256976 7936
rect 131816 7896 131822 7908
rect 256970 7896 256976 7908
rect 257028 7896 257034 7948
rect 77386 7828 77392 7880
rect 77444 7868 77450 7880
rect 218146 7868 218152 7880
rect 77444 7840 218152 7868
rect 77444 7828 77450 7840
rect 218146 7828 218152 7840
rect 218204 7828 218210 7880
rect 73798 7760 73804 7812
rect 73856 7800 73862 7812
rect 215294 7800 215300 7812
rect 73856 7772 215300 7800
rect 73856 7760 73862 7772
rect 215294 7760 215300 7772
rect 215352 7760 215358 7812
rect 343358 7760 343364 7812
rect 343416 7800 343422 7812
rect 409966 7800 409972 7812
rect 343416 7772 409972 7800
rect 343416 7760 343422 7772
rect 409966 7760 409972 7772
rect 410024 7760 410030 7812
rect 38378 7692 38384 7744
rect 38436 7732 38442 7744
rect 180058 7732 180064 7744
rect 38436 7704 180064 7732
rect 38436 7692 38442 7704
rect 180058 7692 180064 7704
rect 180116 7692 180122 7744
rect 181438 7692 181444 7744
rect 181496 7732 181502 7744
rect 292758 7732 292764 7744
rect 181496 7704 292764 7732
rect 181496 7692 181502 7704
rect 292758 7692 292764 7704
rect 292816 7692 292822 7744
rect 304350 7692 304356 7744
rect 304408 7732 304414 7744
rect 380986 7732 380992 7744
rect 304408 7704 380992 7732
rect 304408 7692 304414 7704
rect 380986 7692 380992 7704
rect 381044 7692 381050 7744
rect 70302 7624 70308 7676
rect 70360 7664 70366 7676
rect 212718 7664 212724 7676
rect 70360 7636 212724 7664
rect 70360 7624 70366 7636
rect 212718 7624 212724 7636
rect 212776 7624 212782 7676
rect 298370 7624 298376 7676
rect 298428 7664 298434 7676
rect 376846 7664 376852 7676
rect 298428 7636 376852 7664
rect 298428 7624 298434 7636
rect 376846 7624 376852 7636
rect 376904 7624 376910 7676
rect 66714 7556 66720 7608
rect 66772 7596 66778 7608
rect 209866 7596 209872 7608
rect 66772 7568 209872 7596
rect 66772 7556 66778 7568
rect 209866 7556 209872 7568
rect 209924 7556 209930 7608
rect 292482 7556 292488 7608
rect 292540 7596 292546 7608
rect 371234 7596 371240 7608
rect 292540 7568 371240 7596
rect 292540 7556 292546 7568
rect 371234 7556 371240 7568
rect 371292 7556 371298 7608
rect 377674 7556 377680 7608
rect 377732 7596 377738 7608
rect 434806 7596 434812 7608
rect 377732 7568 434812 7596
rect 377732 7556 377738 7568
rect 434806 7556 434812 7568
rect 434864 7556 434870 7608
rect 174262 7488 174268 7540
rect 174320 7528 174326 7540
rect 287146 7528 287152 7540
rect 174320 7500 287152 7528
rect 174320 7488 174326 7500
rect 287146 7488 287152 7500
rect 287204 7488 287210 7540
rect 184934 7420 184940 7472
rect 184992 7460 184998 7472
rect 295334 7460 295340 7472
rect 184992 7432 295340 7460
rect 184992 7420 184998 7432
rect 295334 7420 295340 7432
rect 295392 7420 295398 7472
rect 188522 7352 188528 7404
rect 188580 7392 188586 7404
rect 298094 7392 298100 7404
rect 188580 7364 298100 7392
rect 188580 7352 188586 7364
rect 298094 7352 298100 7364
rect 298152 7352 298158 7404
rect 192018 7284 192024 7336
rect 192076 7324 192082 7336
rect 300854 7324 300860 7336
rect 192076 7296 300860 7324
rect 192076 7284 192082 7296
rect 300854 7284 300860 7296
rect 300912 7284 300918 7336
rect 195606 7216 195612 7268
rect 195664 7256 195670 7268
rect 303614 7256 303620 7268
rect 195664 7228 303620 7256
rect 195664 7216 195670 7228
rect 303614 7216 303620 7228
rect 303672 7216 303678 7268
rect 199102 7148 199108 7200
rect 199160 7188 199166 7200
rect 305086 7188 305092 7200
rect 199160 7160 305092 7188
rect 199160 7148 199166 7160
rect 305086 7148 305092 7160
rect 305144 7148 305150 7200
rect 202690 7080 202696 7132
rect 202748 7120 202754 7132
rect 307846 7120 307852 7132
rect 202748 7092 307852 7120
rect 202748 7080 202754 7092
rect 307846 7080 307852 7092
rect 307904 7080 307910 7132
rect 206186 7012 206192 7064
rect 206244 7052 206250 7064
rect 310606 7052 310612 7064
rect 206244 7024 310612 7052
rect 206244 7012 206250 7024
rect 310606 7012 310612 7024
rect 310664 7012 310670 7064
rect 63218 6808 63224 6860
rect 63276 6848 63282 6860
rect 207106 6848 207112 6860
rect 63276 6820 207112 6848
rect 63276 6808 63282 6820
rect 207106 6808 207112 6820
rect 207164 6808 207170 6860
rect 215662 6808 215668 6860
rect 215720 6848 215726 6860
rect 317414 6848 317420 6860
rect 215720 6820 317420 6848
rect 215720 6808 215726 6820
rect 317414 6808 317420 6820
rect 317472 6808 317478 6860
rect 59630 6740 59636 6792
rect 59688 6780 59694 6792
rect 205634 6780 205640 6792
rect 59688 6752 205640 6780
rect 59688 6740 59694 6752
rect 205634 6740 205640 6752
rect 205692 6740 205698 6792
rect 212166 6740 212172 6792
rect 212224 6780 212230 6792
rect 314654 6780 314660 6792
rect 212224 6752 314660 6780
rect 212224 6740 212230 6752
rect 314654 6740 314660 6752
rect 314712 6740 314718 6792
rect 56042 6672 56048 6724
rect 56100 6712 56106 6724
rect 202966 6712 202972 6724
rect 56100 6684 202972 6712
rect 56100 6672 56106 6684
rect 202966 6672 202972 6684
rect 203024 6672 203030 6724
rect 208578 6672 208584 6724
rect 208636 6712 208642 6724
rect 311894 6712 311900 6724
rect 208636 6684 311900 6712
rect 208636 6672 208642 6684
rect 311894 6672 311900 6684
rect 311952 6672 311958 6724
rect 52546 6604 52552 6656
rect 52604 6644 52610 6656
rect 200206 6644 200212 6656
rect 52604 6616 200212 6644
rect 52604 6604 52610 6616
rect 200206 6604 200212 6616
rect 200264 6604 200270 6656
rect 205082 6604 205088 6656
rect 205140 6644 205146 6656
rect 309134 6644 309140 6656
rect 205140 6616 309140 6644
rect 205140 6604 205146 6616
rect 309134 6604 309140 6616
rect 309192 6604 309198 6656
rect 48958 6536 48964 6588
rect 49016 6576 49022 6588
rect 197354 6576 197360 6588
rect 49016 6548 197360 6576
rect 49016 6536 49022 6548
rect 197354 6536 197360 6548
rect 197412 6536 197418 6588
rect 201494 6536 201500 6588
rect 201552 6576 201558 6588
rect 307754 6576 307760 6588
rect 201552 6548 307760 6576
rect 201552 6536 201558 6548
rect 307754 6536 307760 6548
rect 307812 6536 307818 6588
rect 44266 6468 44272 6520
rect 44324 6508 44330 6520
rect 194594 6508 194600 6520
rect 44324 6480 194600 6508
rect 44324 6468 44330 6480
rect 194594 6468 194600 6480
rect 194652 6468 194658 6520
rect 197906 6468 197912 6520
rect 197964 6508 197970 6520
rect 304994 6508 305000 6520
rect 197964 6480 305000 6508
rect 197964 6468 197970 6480
rect 304994 6468 305000 6480
rect 305052 6468 305058 6520
rect 40770 6400 40776 6452
rect 40828 6440 40834 6452
rect 191834 6440 191840 6452
rect 40828 6412 191840 6440
rect 40828 6400 40834 6412
rect 191834 6400 191840 6412
rect 191892 6400 191898 6452
rect 194410 6400 194416 6452
rect 194468 6440 194474 6452
rect 302234 6440 302240 6452
rect 194468 6412 302240 6440
rect 194468 6400 194474 6412
rect 302234 6400 302240 6412
rect 302292 6400 302298 6452
rect 345750 6400 345756 6452
rect 345808 6440 345814 6452
rect 411254 6440 411260 6452
rect 345808 6412 411260 6440
rect 345808 6400 345814 6412
rect 411254 6400 411260 6412
rect 411312 6400 411318 6452
rect 37182 6332 37188 6384
rect 37240 6372 37246 6384
rect 189166 6372 189172 6384
rect 37240 6344 189172 6372
rect 37240 6332 37246 6344
rect 189166 6332 189172 6344
rect 189224 6332 189230 6384
rect 190822 6332 190828 6384
rect 190880 6372 190886 6384
rect 299566 6372 299572 6384
rect 190880 6344 299572 6372
rect 190880 6332 190886 6344
rect 299566 6332 299572 6344
rect 299624 6332 299630 6384
rect 339862 6332 339868 6384
rect 339920 6372 339926 6384
rect 407206 6372 407212 6384
rect 339920 6344 407212 6372
rect 339920 6332 339926 6344
rect 407206 6332 407212 6344
rect 407264 6332 407270 6384
rect 33594 6264 33600 6316
rect 33652 6304 33658 6316
rect 186314 6304 186320 6316
rect 33652 6276 186320 6304
rect 33652 6264 33658 6276
rect 186314 6264 186320 6276
rect 186372 6264 186378 6316
rect 187326 6264 187332 6316
rect 187384 6304 187390 6316
rect 296714 6304 296720 6316
rect 187384 6276 296720 6304
rect 187384 6264 187390 6276
rect 296714 6264 296720 6276
rect 296772 6264 296778 6316
rect 335078 6264 335084 6316
rect 335136 6304 335142 6316
rect 403066 6304 403072 6316
rect 335136 6276 403072 6304
rect 335136 6264 335142 6276
rect 403066 6264 403072 6276
rect 403124 6264 403130 6316
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 168374 6236 168380 6248
rect 8812 6208 168380 6236
rect 8812 6196 8818 6208
rect 168374 6196 168380 6208
rect 168432 6196 168438 6248
rect 173158 6196 173164 6248
rect 173216 6236 173222 6248
rect 287054 6236 287060 6248
rect 173216 6208 287060 6236
rect 173216 6196 173222 6208
rect 287054 6196 287060 6208
rect 287112 6196 287118 6248
rect 318518 6196 318524 6248
rect 318576 6236 318582 6248
rect 392026 6236 392032 6248
rect 318576 6208 392032 6236
rect 318576 6196 318582 6208
rect 392026 6196 392032 6208
rect 392084 6196 392090 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 165706 6168 165712 6180
rect 4120 6140 165712 6168
rect 4120 6128 4126 6140
rect 165706 6128 165712 6140
rect 165764 6128 165770 6180
rect 169570 6128 169576 6180
rect 169628 6168 169634 6180
rect 284294 6168 284300 6180
rect 169628 6140 284300 6168
rect 169628 6128 169634 6140
rect 284294 6128 284300 6140
rect 284352 6128 284358 6180
rect 307938 6128 307944 6180
rect 307996 6168 308002 6180
rect 383010 6168 383016 6180
rect 307996 6140 383016 6168
rect 307996 6128 308002 6140
rect 383010 6128 383016 6140
rect 383068 6128 383074 6180
rect 445754 6128 445760 6180
rect 445812 6168 445818 6180
rect 483106 6168 483112 6180
rect 445812 6140 483112 6168
rect 445812 6128 445818 6140
rect 483106 6128 483112 6140
rect 483164 6128 483170 6180
rect 101030 6060 101036 6112
rect 101088 6100 101094 6112
rect 234798 6100 234804 6112
rect 101088 6072 234804 6100
rect 101088 6060 101094 6072
rect 234798 6060 234804 6072
rect 234856 6060 234862 6112
rect 271230 6060 271236 6112
rect 271288 6100 271294 6112
rect 357526 6100 357532 6112
rect 271288 6072 357532 6100
rect 271288 6060 271294 6072
rect 357526 6060 357532 6072
rect 357584 6060 357590 6112
rect 126974 5992 126980 6044
rect 127032 6032 127038 6044
rect 254026 6032 254032 6044
rect 127032 6004 254032 6032
rect 127032 5992 127038 6004
rect 254026 5992 254032 6004
rect 254084 5992 254090 6044
rect 274818 5992 274824 6044
rect 274876 6032 274882 6044
rect 360194 6032 360200 6044
rect 274876 6004 360200 6032
rect 274876 5992 274882 6004
rect 360194 5992 360200 6004
rect 360252 5992 360258 6044
rect 130562 5924 130568 5976
rect 130620 5964 130626 5976
rect 256694 5964 256700 5976
rect 130620 5936 256700 5964
rect 130620 5924 130626 5936
rect 256694 5924 256700 5936
rect 256752 5924 256758 5976
rect 278314 5924 278320 5976
rect 278372 5964 278378 5976
rect 362954 5964 362960 5976
rect 278372 5936 362960 5964
rect 278372 5924 278378 5936
rect 362954 5924 362960 5936
rect 363012 5924 363018 5976
rect 162486 5856 162492 5908
rect 162544 5896 162550 5908
rect 278866 5896 278872 5908
rect 162544 5868 278872 5896
rect 162544 5856 162550 5868
rect 278866 5856 278872 5868
rect 278924 5856 278930 5908
rect 166074 5788 166080 5840
rect 166132 5828 166138 5840
rect 281718 5828 281724 5840
rect 166132 5800 281724 5828
rect 166132 5788 166138 5800
rect 281718 5788 281724 5800
rect 281776 5788 281782 5840
rect 176654 5720 176660 5772
rect 176712 5760 176718 5772
rect 289814 5760 289820 5772
rect 176712 5732 289820 5760
rect 176712 5720 176718 5732
rect 289814 5720 289820 5732
rect 289872 5720 289878 5772
rect 180242 5652 180248 5704
rect 180300 5692 180306 5704
rect 292574 5692 292580 5704
rect 180300 5664 292580 5692
rect 180300 5652 180306 5664
rect 292574 5652 292580 5664
rect 292632 5652 292638 5704
rect 183738 5584 183744 5636
rect 183796 5624 183802 5636
rect 293954 5624 293960 5636
rect 183796 5596 293960 5624
rect 183796 5584 183802 5596
rect 293954 5584 293960 5596
rect 294012 5584 294018 5636
rect 69106 5448 69112 5500
rect 69164 5488 69170 5500
rect 212534 5488 212540 5500
rect 69164 5460 212540 5488
rect 69164 5448 69170 5460
rect 212534 5448 212540 5460
rect 212592 5448 212598 5500
rect 303154 5448 303160 5500
rect 303212 5488 303218 5500
rect 380894 5488 380900 5500
rect 303212 5460 380900 5488
rect 303212 5448 303218 5460
rect 380894 5448 380900 5460
rect 380952 5448 380958 5500
rect 65518 5380 65524 5432
rect 65576 5420 65582 5432
rect 209774 5420 209780 5432
rect 65576 5392 209780 5420
rect 65576 5380 65582 5392
rect 209774 5380 209780 5392
rect 209832 5380 209838 5432
rect 292574 5380 292580 5432
rect 292632 5420 292638 5432
rect 372798 5420 372804 5432
rect 292632 5392 372804 5420
rect 292632 5380 292638 5392
rect 372798 5380 372804 5392
rect 372856 5380 372862 5432
rect 62022 5312 62028 5364
rect 62080 5352 62086 5364
rect 207014 5352 207020 5364
rect 62080 5324 207020 5352
rect 62080 5312 62086 5324
rect 207014 5312 207020 5324
rect 207072 5312 207078 5364
rect 288986 5312 288992 5364
rect 289044 5352 289050 5364
rect 369946 5352 369952 5364
rect 289044 5324 369952 5352
rect 289044 5312 289050 5324
rect 369946 5312 369952 5324
rect 370004 5312 370010 5364
rect 58434 5244 58440 5296
rect 58492 5284 58498 5296
rect 204254 5284 204260 5296
rect 58492 5256 204260 5284
rect 58492 5244 58498 5256
rect 204254 5244 204260 5256
rect 204312 5244 204318 5296
rect 285398 5244 285404 5296
rect 285456 5284 285462 5296
rect 367186 5284 367192 5296
rect 285456 5256 367192 5284
rect 285456 5244 285462 5256
rect 367186 5244 367192 5256
rect 367244 5244 367250 5296
rect 54938 5176 54944 5228
rect 54996 5216 55002 5228
rect 201586 5216 201592 5228
rect 54996 5188 201592 5216
rect 54996 5176 55002 5188
rect 201586 5176 201592 5188
rect 201644 5176 201650 5228
rect 216858 5176 216864 5228
rect 216916 5216 216922 5228
rect 276658 5216 276664 5228
rect 216916 5188 276664 5216
rect 216916 5176 216922 5188
rect 276658 5176 276664 5188
rect 276716 5176 276722 5228
rect 281902 5176 281908 5228
rect 281960 5216 281966 5228
rect 365714 5216 365720 5228
rect 281960 5188 365720 5216
rect 281960 5176 281966 5188
rect 365714 5176 365720 5188
rect 365772 5176 365778 5228
rect 51350 5108 51356 5160
rect 51408 5148 51414 5160
rect 199010 5148 199016 5160
rect 51408 5120 199016 5148
rect 51408 5108 51414 5120
rect 199010 5108 199016 5120
rect 199068 5108 199074 5160
rect 209774 5108 209780 5160
rect 209832 5148 209838 5160
rect 295978 5148 295984 5160
rect 209832 5120 295984 5148
rect 209832 5108 209838 5120
rect 295978 5108 295984 5120
rect 296036 5108 296042 5160
rect 296070 5108 296076 5160
rect 296128 5148 296134 5160
rect 375374 5148 375380 5160
rect 296128 5120 375380 5148
rect 296128 5108 296134 5120
rect 375374 5108 375380 5120
rect 375432 5108 375438 5160
rect 26510 5040 26516 5092
rect 26568 5080 26574 5092
rect 180886 5080 180892 5092
rect 26568 5052 180892 5080
rect 26568 5040 26574 5052
rect 180886 5040 180892 5052
rect 180944 5040 180950 5092
rect 257062 5040 257068 5092
rect 257120 5080 257126 5092
rect 347774 5080 347780 5092
rect 257120 5052 347780 5080
rect 257120 5040 257126 5052
rect 347774 5040 347780 5052
rect 347832 5040 347838 5092
rect 30098 4972 30104 5024
rect 30156 5012 30162 5024
rect 183646 5012 183652 5024
rect 30156 4984 183652 5012
rect 30156 4972 30162 4984
rect 183646 4972 183652 4984
rect 183704 4972 183710 5024
rect 260650 4972 260656 5024
rect 260708 5012 260714 5024
rect 350534 5012 350540 5024
rect 260708 4984 350540 5012
rect 260708 4972 260714 4984
rect 350534 4972 350540 4984
rect 350592 4972 350598 5024
rect 21818 4904 21824 4956
rect 21876 4944 21882 4956
rect 178034 4944 178040 4956
rect 21876 4916 178040 4944
rect 21876 4904 21882 4916
rect 178034 4904 178040 4916
rect 178092 4904 178098 4956
rect 253474 4904 253480 4956
rect 253532 4944 253538 4956
rect 345014 4944 345020 4956
rect 253532 4916 345020 4944
rect 253532 4904 253538 4916
rect 345014 4904 345020 4916
rect 345072 4904 345078 4956
rect 17034 4836 17040 4888
rect 17092 4876 17098 4888
rect 173986 4876 173992 4888
rect 17092 4848 173992 4876
rect 17092 4836 17098 4848
rect 173986 4836 173992 4848
rect 174044 4836 174050 4888
rect 246390 4836 246396 4888
rect 246448 4876 246454 4888
rect 339586 4876 339592 4888
rect 246448 4848 339592 4876
rect 246448 4836 246454 4848
rect 339586 4836 339592 4848
rect 339644 4836 339650 4888
rect 384758 4836 384764 4888
rect 384816 4876 384822 4888
rect 438946 4876 438952 4888
rect 384816 4848 438952 4876
rect 384816 4836 384822 4848
rect 438946 4836 438952 4848
rect 439004 4836 439010 4888
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 171134 4808 171140 4820
rect 12400 4780 171140 4808
rect 12400 4768 12406 4780
rect 171134 4768 171140 4780
rect 171192 4768 171198 4820
rect 242894 4768 242900 4820
rect 242952 4808 242958 4820
rect 337010 4808 337016 4820
rect 242952 4780 337016 4808
rect 242952 4768 242958 4780
rect 337010 4768 337016 4780
rect 337068 4768 337074 4820
rect 370590 4768 370596 4820
rect 370648 4808 370654 4820
rect 429194 4808 429200 4820
rect 370648 4780 429200 4808
rect 370648 4768 370654 4780
rect 429194 4768 429200 4780
rect 429252 4768 429258 4820
rect 72602 4700 72608 4752
rect 72660 4740 72666 4752
rect 214006 4740 214012 4752
rect 72660 4712 214012 4740
rect 72660 4700 72666 4712
rect 214006 4700 214012 4712
rect 214064 4700 214070 4752
rect 299658 4700 299664 4752
rect 299716 4740 299722 4752
rect 378134 4740 378140 4752
rect 299716 4712 378140 4740
rect 299716 4700 299722 4712
rect 378134 4700 378140 4712
rect 378192 4700 378198 4752
rect 79686 4632 79692 4684
rect 79744 4672 79750 4684
rect 219526 4672 219532 4684
rect 79744 4644 219532 4672
rect 79744 4632 79750 4644
rect 219526 4632 219532 4644
rect 219584 4632 219590 4684
rect 306742 4632 306748 4684
rect 306800 4672 306806 4684
rect 383746 4672 383752 4684
rect 306800 4644 383752 4672
rect 306800 4632 306806 4644
rect 383746 4632 383752 4644
rect 383804 4632 383810 4684
rect 76190 4564 76196 4616
rect 76248 4604 76254 4616
rect 216950 4604 216956 4616
rect 76248 4576 216956 4604
rect 76248 4564 76254 4576
rect 216950 4564 216956 4576
rect 217008 4564 217014 4616
rect 310238 4564 310244 4616
rect 310296 4604 310302 4616
rect 385126 4604 385132 4616
rect 310296 4576 385132 4604
rect 310296 4564 310302 4576
rect 385126 4564 385132 4576
rect 385184 4564 385190 4616
rect 86862 4496 86868 4548
rect 86920 4536 86926 4548
rect 224954 4536 224960 4548
rect 86920 4508 224960 4536
rect 86920 4496 86926 4508
rect 224954 4496 224960 4508
rect 225012 4496 225018 4548
rect 317322 4496 317328 4548
rect 317380 4536 317386 4548
rect 390738 4536 390744 4548
rect 317380 4508 390744 4536
rect 317380 4496 317386 4508
rect 390738 4496 390744 4508
rect 390796 4496 390802 4548
rect 83274 4428 83280 4480
rect 83332 4468 83338 4480
rect 222194 4468 222200 4480
rect 83332 4440 222200 4468
rect 83332 4428 83338 4440
rect 222194 4428 222200 4440
rect 222252 4428 222258 4480
rect 313826 4428 313832 4480
rect 313884 4468 313890 4480
rect 387886 4468 387892 4480
rect 313884 4440 387892 4468
rect 313884 4428 313890 4440
rect 387886 4428 387892 4440
rect 387944 4428 387950 4480
rect 90358 4360 90364 4412
rect 90416 4400 90422 4412
rect 227714 4400 227720 4412
rect 90416 4372 227720 4400
rect 90416 4360 90422 4372
rect 227714 4360 227720 4372
rect 227772 4360 227778 4412
rect 320910 4360 320916 4412
rect 320968 4400 320974 4412
rect 393314 4400 393320 4412
rect 320968 4372 393320 4400
rect 320968 4360 320974 4372
rect 393314 4360 393320 4372
rect 393372 4360 393378 4412
rect 93946 4292 93952 4344
rect 94004 4332 94010 4344
rect 229186 4332 229192 4344
rect 94004 4304 229192 4332
rect 94004 4292 94010 4304
rect 229186 4292 229192 4304
rect 229244 4292 229250 4344
rect 327994 4292 328000 4344
rect 328052 4332 328058 4344
rect 398834 4332 398840 4344
rect 328052 4304 398840 4332
rect 328052 4292 328058 4304
rect 398834 4292 398840 4304
rect 398892 4292 398898 4344
rect 97442 4224 97448 4276
rect 97500 4264 97506 4276
rect 231946 4264 231952 4276
rect 97500 4236 231952 4264
rect 97500 4224 97506 4236
rect 231946 4224 231952 4236
rect 232004 4224 232010 4276
rect 324406 4224 324412 4276
rect 324464 4264 324470 4276
rect 396074 4264 396080 4276
rect 324464 4236 396080 4264
rect 324464 4224 324470 4236
rect 396074 4224 396080 4236
rect 396132 4224 396138 4276
rect 402440 4168 403112 4196
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 18598 4128 18604 4140
rect 14792 4100 18604 4128
rect 14792 4088 14798 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 33778 4128 33784 4140
rect 18800 4100 33784 4128
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 18800 4060 18828 4100
rect 33778 4088 33784 4100
rect 33836 4088 33842 4140
rect 36538 4128 36544 4140
rect 33888 4100 36544 4128
rect 18288 4032 18828 4060
rect 18288 4020 18294 4032
rect 25314 4020 25320 4072
rect 25372 4060 25378 4072
rect 29638 4060 29644 4072
rect 25372 4032 29644 4060
rect 25372 4020 25378 4032
rect 29638 4020 29644 4032
rect 29696 4020 29702 4072
rect 32398 4020 32404 4072
rect 32456 4060 32462 4072
rect 33888 4060 33916 4100
rect 36538 4088 36544 4100
rect 36596 4088 36602 4140
rect 57238 4128 57244 4140
rect 40696 4100 57244 4128
rect 32456 4032 33916 4060
rect 32456 4020 32462 4032
rect 34790 4020 34796 4072
rect 34848 4060 34854 4072
rect 40696 4060 40724 4100
rect 57238 4088 57244 4100
rect 57296 4088 57302 4140
rect 67910 4088 67916 4140
rect 67968 4128 67974 4140
rect 195238 4128 195244 4140
rect 67968 4100 195244 4128
rect 67968 4088 67974 4100
rect 195238 4088 195244 4100
rect 195296 4088 195302 4140
rect 214466 4088 214472 4140
rect 214524 4128 214530 4140
rect 228177 4131 228235 4137
rect 228177 4128 228189 4131
rect 214524 4100 228189 4128
rect 214524 4088 214530 4100
rect 228177 4097 228189 4100
rect 228223 4097 228235 4131
rect 228177 4091 228235 4097
rect 229830 4088 229836 4140
rect 229888 4128 229894 4140
rect 233970 4128 233976 4140
rect 229888 4100 233976 4128
rect 229888 4088 229894 4100
rect 233970 4088 233976 4100
rect 234028 4088 234034 4140
rect 237006 4088 237012 4140
rect 237064 4128 237070 4140
rect 239217 4131 239275 4137
rect 237064 4100 239168 4128
rect 237064 4088 237070 4100
rect 34848 4032 40724 4060
rect 40773 4063 40831 4069
rect 34848 4020 34854 4032
rect 40773 4029 40785 4063
rect 40819 4060 40831 4063
rect 54478 4060 54484 4072
rect 40819 4032 54484 4060
rect 40819 4029 40831 4032
rect 40773 4023 40831 4029
rect 54478 4020 54484 4032
rect 54536 4020 54542 4072
rect 60826 4020 60832 4072
rect 60884 4060 60890 4072
rect 192478 4060 192484 4072
rect 60884 4032 192484 4060
rect 60884 4020 60890 4032
rect 192478 4020 192484 4032
rect 192536 4020 192542 4072
rect 207382 4020 207388 4072
rect 207440 4060 207446 4072
rect 239033 4063 239091 4069
rect 239033 4060 239045 4063
rect 207440 4032 239045 4060
rect 207440 4020 207446 4032
rect 239033 4029 239045 4032
rect 239079 4029 239091 4063
rect 239140 4060 239168 4100
rect 239217 4097 239229 4131
rect 239263 4128 239275 4131
rect 313918 4128 313924 4140
rect 239263 4100 313924 4128
rect 239263 4097 239275 4100
rect 239217 4091 239275 4097
rect 313918 4088 313924 4100
rect 313976 4088 313982 4140
rect 316218 4088 316224 4140
rect 316276 4128 316282 4140
rect 389818 4128 389824 4140
rect 316276 4100 389824 4128
rect 316276 4088 316282 4100
rect 389818 4088 389824 4100
rect 389876 4088 389882 4140
rect 393038 4088 393044 4140
rect 393096 4128 393102 4140
rect 393958 4128 393964 4140
rect 393096 4100 393964 4128
rect 393096 4088 393102 4100
rect 393958 4088 393964 4100
rect 394016 4088 394022 4140
rect 396721 4131 396779 4137
rect 396721 4097 396733 4131
rect 396767 4128 396779 4131
rect 400214 4128 400220 4140
rect 396767 4100 400220 4128
rect 396767 4097 396779 4100
rect 396721 4091 396779 4097
rect 400214 4088 400220 4100
rect 400272 4088 400278 4140
rect 401318 4088 401324 4140
rect 401376 4128 401382 4140
rect 402440 4128 402468 4168
rect 401376 4100 402468 4128
rect 401376 4088 401382 4100
rect 402514 4088 402520 4140
rect 402572 4128 402578 4140
rect 402974 4128 402980 4140
rect 402572 4100 402980 4128
rect 402572 4088 402578 4100
rect 402974 4088 402980 4100
rect 403032 4088 403038 4140
rect 403084 4128 403112 4168
rect 451274 4128 451280 4140
rect 403084 4100 451280 4128
rect 451274 4088 451280 4100
rect 451332 4088 451338 4140
rect 456886 4088 456892 4140
rect 456944 4128 456950 4140
rect 461578 4128 461584 4140
rect 456944 4100 461584 4128
rect 456944 4088 456950 4100
rect 461578 4088 461584 4100
rect 461636 4088 461642 4140
rect 465721 4131 465779 4137
rect 465721 4097 465733 4131
rect 465767 4128 465779 4131
rect 473998 4128 474004 4140
rect 465767 4100 474004 4128
rect 465767 4097 465779 4100
rect 465721 4091 465779 4097
rect 473998 4088 474004 4100
rect 474056 4088 474062 4140
rect 497090 4088 497096 4140
rect 497148 4128 497154 4140
rect 501598 4128 501604 4140
rect 497148 4100 501604 4128
rect 497148 4088 497154 4100
rect 501598 4088 501604 4100
rect 501656 4088 501662 4140
rect 556154 4088 556160 4140
rect 556212 4128 556218 4140
rect 558270 4128 558276 4140
rect 556212 4100 558276 4128
rect 556212 4088 556218 4100
rect 558270 4088 558276 4100
rect 558328 4088 558334 4140
rect 240778 4060 240784 4072
rect 239140 4032 240784 4060
rect 239033 4023 239091 4029
rect 240778 4020 240784 4032
rect 240836 4020 240842 4072
rect 247586 4020 247592 4072
rect 247644 4060 247650 4072
rect 273898 4060 273904 4072
rect 247644 4032 273904 4060
rect 247644 4020 247650 4032
rect 273898 4020 273904 4032
rect 273956 4020 273962 4072
rect 280706 4020 280712 4072
rect 280764 4060 280770 4072
rect 286413 4063 286471 4069
rect 286413 4060 286425 4063
rect 280764 4032 286425 4060
rect 280764 4020 280770 4032
rect 286413 4029 286425 4032
rect 286459 4029 286471 4063
rect 286413 4023 286471 4029
rect 287790 4020 287796 4072
rect 287848 4060 287854 4072
rect 287848 4032 293356 4060
rect 287848 4020 287854 4032
rect 1670 3952 1676 4004
rect 1728 3992 1734 4004
rect 22738 3992 22744 4004
rect 1728 3964 22744 3992
rect 1728 3952 1734 3964
rect 22738 3952 22744 3964
rect 22796 3952 22802 4004
rect 27706 3952 27712 4004
rect 27764 3992 27770 4004
rect 51718 3992 51724 4004
rect 27764 3964 51724 3992
rect 27764 3952 27770 3964
rect 51718 3952 51724 3964
rect 51776 3952 51782 4004
rect 53742 3952 53748 4004
rect 53800 3992 53806 4004
rect 191098 3992 191104 4004
rect 53800 3964 191104 3992
rect 53800 3952 53806 3964
rect 191098 3952 191104 3964
rect 191156 3952 191162 4004
rect 210970 3952 210976 4004
rect 211028 3992 211034 4004
rect 250438 3992 250444 4004
rect 211028 3964 250444 3992
rect 211028 3952 211034 3964
rect 250438 3952 250444 3964
rect 250496 3952 250502 4004
rect 258166 3952 258172 4004
rect 258224 3992 258230 4004
rect 258810 3992 258816 4004
rect 258224 3964 258816 3992
rect 258224 3952 258230 3964
rect 258810 3952 258816 3964
rect 258868 3952 258874 4004
rect 265342 3952 265348 4004
rect 265400 3992 265406 4004
rect 268378 3992 268384 4004
rect 265400 3964 268384 3992
rect 265400 3952 265406 3964
rect 268378 3952 268384 3964
rect 268436 3952 268442 4004
rect 272426 3952 272432 4004
rect 272484 3992 272490 4004
rect 282178 3992 282184 4004
rect 272484 3964 282184 3992
rect 272484 3952 272490 3964
rect 282178 3952 282184 3964
rect 282236 3952 282242 4004
rect 283098 3952 283104 4004
rect 283156 3992 283162 4004
rect 291286 3992 291292 4004
rect 283156 3964 291292 3992
rect 283156 3952 283162 3964
rect 291286 3952 291292 3964
rect 291344 3952 291350 4004
rect 291378 3952 291384 4004
rect 291436 3992 291442 4004
rect 293218 3992 293224 4004
rect 291436 3964 293224 3992
rect 291436 3952 291442 3964
rect 293218 3952 293224 3964
rect 293276 3952 293282 4004
rect 293328 3992 293356 4032
rect 294874 4020 294880 4072
rect 294932 4060 294938 4072
rect 373994 4060 374000 4072
rect 294932 4032 374000 4060
rect 294932 4020 294938 4032
rect 373994 4020 374000 4032
rect 374052 4020 374058 4072
rect 383562 4020 383568 4072
rect 383620 4060 383626 4072
rect 384298 4060 384304 4072
rect 383620 4032 384304 4060
rect 383620 4020 383626 4032
rect 384298 4020 384304 4032
rect 384356 4020 384362 4072
rect 385954 4020 385960 4072
rect 386012 4060 386018 4072
rect 388438 4060 388444 4072
rect 386012 4032 388444 4060
rect 386012 4020 386018 4032
rect 388438 4020 388444 4032
rect 388496 4020 388502 4072
rect 389450 4020 389456 4072
rect 389508 4060 389514 4072
rect 389508 4032 437796 4060
rect 389508 4020 389514 4032
rect 369854 3992 369860 4004
rect 293328 3964 369860 3992
rect 369854 3952 369860 3964
rect 369912 3952 369918 4004
rect 382366 3952 382372 4004
rect 382424 3992 382430 4004
rect 437658 3992 437664 4004
rect 382424 3964 437664 3992
rect 382424 3952 382430 3964
rect 437658 3952 437664 3964
rect 437716 3952 437722 4004
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 39298 3924 39304 3936
rect 13596 3896 39304 3924
rect 13596 3884 13602 3896
rect 39298 3884 39304 3896
rect 39356 3884 39362 3936
rect 43070 3884 43076 3936
rect 43128 3924 43134 3936
rect 193214 3924 193220 3936
rect 43128 3896 193220 3924
rect 43128 3884 43134 3896
rect 193214 3884 193220 3896
rect 193272 3884 193278 3936
rect 218054 3884 218060 3936
rect 218112 3924 218118 3936
rect 262858 3924 262864 3936
rect 218112 3896 262864 3924
rect 218112 3884 218118 3896
rect 262858 3884 262864 3896
rect 262916 3884 262922 3936
rect 266538 3884 266544 3936
rect 266596 3924 266602 3936
rect 349798 3924 349804 3936
rect 266596 3896 349804 3924
rect 266596 3884 266602 3896
rect 349798 3884 349804 3896
rect 349856 3884 349862 3936
rect 352834 3884 352840 3936
rect 352892 3924 352898 3936
rect 353938 3924 353944 3936
rect 352892 3896 353944 3924
rect 352892 3884 352898 3896
rect 353938 3884 353944 3896
rect 353996 3884 354002 3936
rect 356330 3884 356336 3936
rect 356388 3924 356394 3936
rect 357342 3924 357348 3936
rect 356388 3896 357348 3924
rect 356388 3884 356394 3896
rect 357342 3884 357348 3896
rect 357400 3884 357406 3936
rect 357526 3884 357532 3936
rect 357584 3924 357590 3936
rect 358722 3924 358728 3936
rect 357584 3896 358728 3924
rect 357584 3884 357590 3896
rect 358722 3884 358728 3896
rect 358780 3884 358786 3936
rect 420914 3924 420920 3936
rect 373966 3896 420920 3924
rect 7650 3816 7656 3868
rect 7708 3856 7714 3868
rect 32306 3856 32312 3868
rect 7708 3828 32312 3856
rect 7708 3816 7714 3828
rect 32306 3816 32312 3828
rect 32364 3816 32370 3868
rect 35986 3816 35992 3868
rect 36044 3856 36050 3868
rect 187694 3856 187700 3868
rect 36044 3828 187700 3856
rect 36044 3816 36050 3828
rect 187694 3816 187700 3828
rect 187752 3816 187758 3868
rect 203886 3816 203892 3868
rect 203944 3856 203950 3868
rect 252002 3856 252008 3868
rect 203944 3828 252008 3856
rect 203944 3816 203950 3828
rect 252002 3816 252008 3828
rect 252060 3816 252066 3868
rect 254670 3816 254676 3868
rect 254728 3856 254734 3868
rect 254728 3828 258074 3856
rect 254728 3816 254734 3828
rect 2866 3748 2872 3800
rect 2924 3788 2930 3800
rect 25498 3788 25504 3800
rect 2924 3760 25504 3788
rect 2924 3748 2930 3760
rect 25498 3748 25504 3760
rect 25556 3748 25562 3800
rect 28902 3748 28908 3800
rect 28960 3788 28966 3800
rect 183554 3788 183560 3800
rect 28960 3760 183560 3788
rect 28960 3748 28966 3760
rect 183554 3748 183560 3760
rect 183612 3748 183618 3800
rect 196802 3748 196808 3800
rect 196860 3788 196866 3800
rect 255958 3788 255964 3800
rect 196860 3760 255964 3788
rect 196860 3748 196866 3760
rect 255958 3748 255964 3760
rect 256016 3748 256022 3800
rect 258046 3788 258074 3828
rect 261754 3816 261760 3868
rect 261812 3856 261818 3868
rect 278038 3856 278044 3868
rect 261812 3828 278044 3856
rect 261812 3816 261818 3828
rect 278038 3816 278044 3828
rect 278096 3816 278102 3868
rect 279510 3816 279516 3868
rect 279568 3856 279574 3868
rect 286318 3856 286324 3868
rect 279568 3828 286324 3856
rect 279568 3816 279574 3828
rect 286318 3816 286324 3828
rect 286376 3816 286382 3868
rect 286413 3859 286471 3865
rect 286413 3825 286425 3859
rect 286459 3856 286471 3859
rect 286459 3828 356836 3856
rect 286459 3825 286471 3828
rect 286413 3819 286471 3825
rect 269114 3788 269120 3800
rect 258046 3760 269120 3788
rect 269114 3748 269120 3760
rect 269172 3748 269178 3800
rect 273622 3748 273628 3800
rect 273680 3788 273686 3800
rect 354677 3791 354735 3797
rect 354677 3788 354689 3791
rect 273680 3760 354689 3788
rect 273680 3748 273686 3760
rect 354677 3757 354689 3760
rect 354723 3757 354735 3791
rect 354677 3751 354735 3757
rect 355226 3748 355232 3800
rect 355284 3788 355290 3800
rect 356698 3788 356704 3800
rect 355284 3760 356704 3788
rect 355284 3748 355290 3760
rect 356698 3748 356704 3760
rect 356756 3748 356762 3800
rect 356808 3788 356836 3828
rect 358630 3816 358636 3868
rect 358688 3856 358694 3868
rect 373966 3856 373994 3896
rect 420914 3884 420920 3896
rect 420972 3884 420978 3936
rect 421009 3927 421067 3933
rect 421009 3893 421021 3927
rect 421055 3924 421067 3927
rect 424318 3924 424324 3936
rect 421055 3896 424324 3924
rect 421055 3893 421067 3896
rect 421009 3887 421067 3893
rect 424318 3884 424324 3896
rect 424376 3884 424382 3936
rect 424873 3927 424931 3933
rect 424873 3893 424885 3927
rect 424919 3924 424931 3927
rect 431218 3924 431224 3936
rect 424919 3896 431224 3924
rect 424919 3893 424931 3896
rect 424873 3887 424931 3893
rect 431218 3884 431224 3896
rect 431276 3884 431282 3936
rect 358688 3828 373994 3856
rect 358688 3816 358694 3828
rect 375190 3816 375196 3868
rect 375248 3856 375254 3868
rect 431954 3856 431960 3868
rect 375248 3828 431960 3856
rect 375248 3816 375254 3828
rect 431954 3816 431960 3828
rect 432012 3816 432018 3868
rect 437768 3856 437796 4032
rect 446214 4020 446220 4072
rect 446272 4060 446278 4072
rect 460198 4060 460204 4072
rect 446272 4032 460204 4060
rect 446272 4020 446278 4032
rect 460198 4020 460204 4032
rect 460256 4020 460262 4072
rect 462774 4020 462780 4072
rect 462832 4060 462838 4072
rect 486326 4060 486332 4072
rect 462832 4032 486332 4060
rect 462832 4020 462838 4032
rect 486326 4020 486332 4032
rect 486384 4020 486390 4072
rect 440326 3952 440332 4004
rect 440384 3992 440390 4004
rect 447045 3995 447103 4001
rect 447045 3992 447057 3995
rect 440384 3964 447057 3992
rect 440384 3952 440390 3964
rect 447045 3961 447057 3964
rect 447091 3961 447103 3995
rect 447045 3955 447103 3961
rect 447152 3964 451274 3992
rect 437845 3927 437903 3933
rect 437845 3893 437857 3927
rect 437891 3924 437903 3927
rect 447152 3924 447180 3964
rect 437891 3896 447180 3924
rect 451246 3924 451274 3964
rect 459186 3952 459192 4004
rect 459244 3992 459250 4004
rect 485038 3992 485044 4004
rect 459244 3964 485044 3992
rect 459244 3952 459250 3964
rect 485038 3952 485044 3964
rect 485096 3952 485102 4004
rect 563238 3952 563244 4004
rect 563296 3992 563302 4004
rect 568574 3992 568580 4004
rect 563296 3964 568580 3992
rect 563296 3952 563302 3964
rect 568574 3952 568580 3964
rect 568632 3952 568638 4004
rect 467098 3924 467104 3936
rect 451246 3896 467104 3924
rect 437891 3893 437903 3896
rect 437845 3887 437903 3893
rect 467098 3884 467104 3896
rect 467156 3884 467162 3936
rect 468662 3884 468668 3936
rect 468720 3924 468726 3936
rect 476758 3924 476764 3936
rect 468720 3896 476764 3924
rect 468720 3884 468726 3896
rect 476758 3884 476764 3896
rect 476816 3884 476822 3936
rect 479334 3884 479340 3936
rect 479392 3924 479398 3936
rect 480898 3924 480904 3936
rect 479392 3896 480904 3924
rect 479392 3884 479398 3896
rect 480898 3884 480904 3896
rect 480956 3884 480962 3936
rect 501509 3927 501567 3933
rect 501509 3893 501521 3927
rect 501555 3924 501567 3927
rect 508498 3924 508504 3936
rect 501555 3896 508504 3924
rect 501555 3893 501567 3896
rect 501509 3887 501567 3893
rect 508498 3884 508504 3896
rect 508556 3884 508562 3936
rect 443086 3856 443092 3868
rect 437768 3828 443092 3856
rect 443086 3816 443092 3828
rect 443144 3816 443150 3868
rect 443733 3859 443791 3865
rect 443733 3825 443745 3859
rect 443779 3856 443791 3859
rect 447134 3856 447140 3868
rect 443779 3828 447140 3856
rect 443779 3825 443791 3828
rect 443733 3819 443791 3825
rect 447134 3816 447140 3828
rect 447192 3816 447198 3868
rect 447229 3859 447287 3865
rect 447229 3825 447241 3859
rect 447275 3856 447287 3859
rect 469858 3856 469864 3868
rect 447275 3828 469864 3856
rect 447275 3825 447287 3828
rect 447229 3819 447287 3825
rect 469858 3816 469864 3828
rect 469916 3816 469922 3868
rect 504174 3816 504180 3868
rect 504232 3856 504238 3868
rect 512638 3856 512644 3868
rect 504232 3828 512644 3856
rect 504232 3816 504238 3828
rect 512638 3816 512644 3828
rect 512696 3816 512702 3868
rect 363598 3788 363604 3800
rect 356808 3760 363604 3788
rect 363598 3748 363604 3760
rect 363656 3748 363662 3800
rect 368198 3748 368204 3800
rect 368256 3788 368262 3800
rect 427906 3788 427912 3800
rect 368256 3760 427912 3788
rect 368256 3748 368262 3760
rect 427906 3748 427912 3760
rect 427964 3748 427970 3800
rect 433153 3791 433211 3797
rect 433153 3757 433165 3791
rect 433199 3788 433211 3791
rect 437661 3791 437719 3797
rect 437661 3788 437673 3791
rect 433199 3760 437673 3788
rect 433199 3757 433211 3760
rect 433153 3751 433211 3757
rect 437661 3757 437673 3760
rect 437707 3757 437719 3791
rect 437661 3751 437719 3757
rect 437753 3791 437811 3797
rect 437753 3757 437765 3791
rect 437799 3788 437811 3791
rect 468478 3788 468484 3800
rect 437799 3760 468484 3788
rect 437799 3757 437811 3760
rect 437753 3751 437811 3757
rect 468478 3748 468484 3760
rect 468536 3748 468542 3800
rect 493502 3748 493508 3800
rect 493560 3788 493566 3800
rect 504358 3788 504364 3800
rect 493560 3760 504364 3788
rect 493560 3748 493566 3760
rect 504358 3748 504364 3760
rect 504416 3748 504422 3800
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 176746 3720 176752 3732
rect 19484 3692 176752 3720
rect 19484 3680 19490 3692
rect 176746 3680 176752 3692
rect 176804 3680 176810 3732
rect 189718 3680 189724 3732
rect 189776 3720 189782 3732
rect 253198 3720 253204 3732
rect 189776 3692 253204 3720
rect 189776 3680 189782 3692
rect 253198 3680 253204 3692
rect 253256 3680 253262 3732
rect 259454 3680 259460 3732
rect 259512 3720 259518 3732
rect 349154 3720 349160 3732
rect 259512 3692 349160 3720
rect 259512 3680 259518 3692
rect 349154 3680 349160 3692
rect 349212 3680 349218 3732
rect 354030 3680 354036 3732
rect 354088 3720 354094 3732
rect 416774 3720 416780 3732
rect 354088 3692 416780 3720
rect 354088 3680 354094 3692
rect 416774 3680 416780 3692
rect 416832 3680 416838 3732
rect 420178 3680 420184 3732
rect 420236 3720 420242 3732
rect 421009 3723 421067 3729
rect 421009 3720 421021 3723
rect 420236 3692 421021 3720
rect 420236 3680 420242 3692
rect 421009 3689 421021 3692
rect 421055 3689 421067 3723
rect 421009 3683 421067 3689
rect 421374 3680 421380 3732
rect 421432 3720 421438 3732
rect 464430 3720 464436 3732
rect 421432 3692 464436 3720
rect 421432 3680 421438 3692
rect 464430 3680 464436 3692
rect 464488 3680 464494 3732
rect 473446 3680 473452 3732
rect 473504 3720 473510 3732
rect 493410 3720 493416 3732
rect 473504 3692 493416 3720
rect 473504 3680 473510 3692
rect 493410 3680 493416 3692
rect 493468 3680 493474 3732
rect 498194 3680 498200 3732
rect 498252 3720 498258 3732
rect 501509 3723 501567 3729
rect 501509 3720 501521 3723
rect 498252 3692 501521 3720
rect 498252 3680 498258 3692
rect 501509 3689 501521 3692
rect 501555 3689 501567 3723
rect 501509 3683 501567 3689
rect 501601 3723 501659 3729
rect 501601 3689 501613 3723
rect 501647 3720 501659 3723
rect 503714 3720 503720 3732
rect 501647 3692 503720 3720
rect 501647 3689 501659 3692
rect 501601 3683 501659 3689
rect 503714 3680 503720 3692
rect 503772 3680 503778 3732
rect 539594 3680 539600 3732
rect 539652 3720 539658 3732
rect 550910 3720 550916 3732
rect 539652 3692 550916 3720
rect 539652 3680 539658 3692
rect 550910 3680 550916 3692
rect 550968 3680 550974 3732
rect 566 3612 572 3664
rect 624 3652 630 3664
rect 14458 3652 14464 3664
rect 624 3624 14464 3652
rect 624 3612 630 3624
rect 14458 3612 14464 3624
rect 14516 3612 14522 3664
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 176930 3652 176936 3664
rect 20680 3624 176936 3652
rect 20680 3612 20686 3624
rect 176930 3612 176936 3624
rect 176988 3612 176994 3664
rect 200298 3612 200304 3664
rect 200356 3652 200362 3664
rect 238941 3655 238999 3661
rect 238941 3652 238953 3655
rect 200356 3624 238953 3652
rect 200356 3612 200362 3624
rect 238941 3621 238953 3624
rect 238987 3621 238999 3655
rect 238941 3615 238999 3621
rect 239033 3655 239091 3661
rect 239033 3621 239045 3655
rect 239079 3652 239091 3655
rect 246298 3652 246304 3664
rect 239079 3624 246304 3652
rect 239079 3621 239091 3624
rect 239033 3615 239091 3621
rect 246298 3612 246304 3624
rect 246356 3612 246362 3664
rect 248782 3612 248788 3664
rect 248840 3652 248846 3664
rect 249702 3652 249708 3664
rect 248840 3624 249708 3652
rect 248840 3612 248846 3624
rect 249702 3612 249708 3624
rect 249760 3612 249766 3664
rect 252370 3612 252376 3664
rect 252428 3652 252434 3664
rect 342898 3652 342904 3664
rect 252428 3624 342904 3652
rect 252428 3612 252434 3624
rect 342898 3612 342904 3624
rect 342956 3612 342962 3664
rect 351638 3612 351644 3664
rect 351696 3652 351702 3664
rect 415394 3652 415400 3664
rect 351696 3624 415400 3652
rect 351696 3612 351702 3624
rect 415394 3612 415400 3624
rect 415452 3612 415458 3664
rect 415489 3655 415547 3661
rect 415489 3621 415501 3655
rect 415535 3652 415547 3655
rect 421558 3652 421564 3664
rect 415535 3624 421564 3652
rect 415535 3621 415547 3624
rect 415489 3615 415547 3621
rect 421558 3612 421564 3624
rect 421616 3612 421622 3664
rect 423677 3655 423735 3661
rect 423677 3621 423689 3655
rect 423723 3652 423735 3655
rect 424873 3655 424931 3661
rect 424873 3652 424885 3655
rect 423723 3624 424885 3652
rect 423723 3621 423735 3624
rect 423677 3615 423735 3621
rect 424873 3621 424885 3624
rect 424919 3621 424931 3655
rect 424873 3615 424931 3621
rect 424962 3612 424968 3664
rect 425020 3652 425026 3664
rect 467834 3652 467840 3664
rect 425020 3624 467840 3652
rect 425020 3612 425026 3624
rect 467834 3612 467840 3624
rect 467892 3612 467898 3664
rect 471517 3655 471575 3661
rect 471517 3621 471529 3655
rect 471563 3652 471575 3655
rect 475378 3652 475384 3664
rect 471563 3624 475384 3652
rect 471563 3621 471575 3624
rect 471517 3615 471575 3621
rect 475378 3612 475384 3624
rect 475436 3612 475442 3664
rect 476942 3612 476948 3664
rect 477000 3652 477006 3664
rect 502886 3652 502892 3664
rect 477000 3624 502892 3652
rect 477000 3612 477006 3624
rect 502886 3612 502892 3624
rect 502944 3612 502950 3664
rect 510614 3652 510620 3664
rect 504376 3624 510620 3652
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 169754 3584 169760 3596
rect 11204 3556 169760 3584
rect 11204 3544 11210 3556
rect 169754 3544 169760 3556
rect 169812 3544 169818 3596
rect 182542 3544 182548 3596
rect 182600 3584 182606 3596
rect 209038 3584 209044 3596
rect 182600 3556 209044 3584
rect 182600 3544 182606 3556
rect 209038 3544 209044 3556
rect 209096 3544 209102 3596
rect 213362 3544 213368 3596
rect 213420 3584 213426 3596
rect 215938 3584 215944 3596
rect 213420 3556 215944 3584
rect 213420 3544 213426 3556
rect 215938 3544 215944 3556
rect 215996 3544 216002 3596
rect 221550 3544 221556 3596
rect 221608 3584 221614 3596
rect 224218 3584 224224 3596
rect 221608 3556 224224 3584
rect 221608 3544 221614 3556
rect 224218 3544 224224 3556
rect 224276 3544 224282 3596
rect 225138 3544 225144 3596
rect 225196 3584 225202 3596
rect 228634 3584 228640 3596
rect 225196 3556 228640 3584
rect 225196 3544 225202 3556
rect 228634 3544 228640 3556
rect 228692 3544 228698 3596
rect 228726 3544 228732 3596
rect 228784 3584 228790 3596
rect 230934 3584 230940 3596
rect 228784 3556 230940 3584
rect 228784 3544 228790 3556
rect 230934 3544 230940 3556
rect 230992 3544 230998 3596
rect 231026 3544 231032 3596
rect 231084 3584 231090 3596
rect 322014 3584 322020 3596
rect 231084 3556 322020 3584
rect 231084 3544 231090 3556
rect 322014 3544 322020 3556
rect 322072 3544 322078 3596
rect 322106 3544 322112 3596
rect 322164 3584 322170 3596
rect 324958 3584 324964 3596
rect 322164 3556 324964 3584
rect 322164 3544 322170 3556
rect 324958 3544 324964 3556
rect 325016 3544 325022 3596
rect 325053 3587 325111 3593
rect 325053 3553 325065 3587
rect 325099 3584 325111 3587
rect 394694 3584 394700 3596
rect 325099 3556 394700 3584
rect 325099 3553 325111 3556
rect 325053 3547 325111 3553
rect 394694 3544 394700 3556
rect 394752 3544 394758 3596
rect 395338 3544 395344 3596
rect 395396 3584 395402 3596
rect 396718 3584 396724 3596
rect 395396 3556 396724 3584
rect 395396 3544 395402 3556
rect 396718 3544 396724 3556
rect 396776 3544 396782 3596
rect 397730 3544 397736 3596
rect 397788 3584 397794 3596
rect 399478 3584 399484 3596
rect 397788 3556 399484 3584
rect 397788 3544 397794 3556
rect 399478 3544 399484 3556
rect 399536 3544 399542 3596
rect 399573 3587 399631 3593
rect 399573 3553 399585 3587
rect 399619 3584 399631 3587
rect 443733 3587 443791 3593
rect 443733 3584 443745 3587
rect 399619 3556 443745 3584
rect 399619 3553 399631 3556
rect 399573 3547 399631 3553
rect 443733 3553 443745 3556
rect 443779 3553 443791 3587
rect 443733 3547 443791 3553
rect 443822 3544 443828 3596
rect 443880 3584 443886 3596
rect 444282 3584 444288 3596
rect 443880 3556 444288 3584
rect 443880 3544 443886 3556
rect 444282 3544 444288 3556
rect 444340 3544 444346 3596
rect 448606 3544 448612 3596
rect 448664 3584 448670 3596
rect 450538 3584 450544 3596
rect 448664 3556 450544 3584
rect 448664 3544 448670 3556
rect 450538 3544 450544 3556
rect 450596 3544 450602 3596
rect 450633 3587 450691 3593
rect 450633 3553 450645 3587
rect 450679 3584 450691 3587
rect 472618 3584 472624 3596
rect 450679 3556 472624 3584
rect 450679 3553 450691 3556
rect 450633 3547 450691 3553
rect 472618 3544 472624 3556
rect 472676 3544 472682 3596
rect 474550 3544 474556 3596
rect 474608 3584 474614 3596
rect 474608 3556 480254 3584
rect 474608 3544 474614 3556
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 164789 3519 164847 3525
rect 164789 3516 164801 3519
rect 10008 3488 164801 3516
rect 10008 3476 10014 3488
rect 164789 3485 164801 3488
rect 164835 3485 164847 3519
rect 164789 3479 164847 3485
rect 164878 3476 164884 3528
rect 164936 3516 164942 3528
rect 165522 3516 165528 3528
rect 164936 3488 165528 3516
rect 164936 3476 164942 3488
rect 165522 3476 165528 3488
rect 165580 3476 165586 3528
rect 168374 3476 168380 3528
rect 168432 3516 168438 3528
rect 169662 3516 169668 3528
rect 168432 3488 169668 3516
rect 168432 3476 168438 3488
rect 169662 3476 169668 3488
rect 169720 3476 169726 3528
rect 175458 3476 175464 3528
rect 175516 3516 175522 3528
rect 176562 3516 176568 3528
rect 175516 3488 176568 3516
rect 175516 3476 175522 3488
rect 176562 3476 176568 3488
rect 176620 3476 176626 3528
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 193272 3488 222700 3516
rect 193272 3476 193278 3488
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 165798 3448 165804 3460
rect 5316 3420 165804 3448
rect 5316 3408 5322 3420
rect 165798 3408 165804 3420
rect 165856 3408 165862 3460
rect 186130 3408 186136 3460
rect 186188 3448 186194 3460
rect 222672 3448 222700 3488
rect 222746 3476 222752 3528
rect 222804 3516 222810 3528
rect 223482 3516 223488 3528
rect 222804 3488 223488 3516
rect 222804 3476 222810 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 224862 3516 224868 3528
rect 224000 3488 224868 3516
rect 224000 3476 224006 3488
rect 224862 3476 224868 3488
rect 224920 3476 224926 3528
rect 228177 3519 228235 3525
rect 228177 3485 228189 3519
rect 228223 3516 228235 3519
rect 234062 3516 234068 3528
rect 228223 3488 234068 3516
rect 228223 3485 228235 3488
rect 228177 3479 228235 3485
rect 234062 3476 234068 3488
rect 234120 3476 234126 3528
rect 234614 3476 234620 3528
rect 234672 3516 234678 3528
rect 239217 3519 239275 3525
rect 239217 3516 239229 3519
rect 234672 3488 239229 3516
rect 234672 3476 234678 3488
rect 239217 3485 239229 3488
rect 239263 3485 239275 3519
rect 239217 3479 239275 3485
rect 239306 3476 239312 3528
rect 239364 3516 239370 3528
rect 240134 3516 240140 3528
rect 239364 3488 240140 3516
rect 239364 3476 239370 3488
rect 240134 3476 240140 3488
rect 240192 3476 240198 3528
rect 241698 3476 241704 3528
rect 241756 3516 241762 3528
rect 242802 3516 242808 3528
rect 241756 3488 242808 3516
rect 241756 3476 241762 3488
rect 242802 3476 242808 3488
rect 242860 3476 242866 3528
rect 245194 3476 245200 3528
rect 245252 3516 245258 3528
rect 338298 3516 338304 3528
rect 245252 3488 338304 3516
rect 245252 3476 245258 3488
rect 338298 3476 338304 3488
rect 338356 3476 338362 3528
rect 338666 3476 338672 3528
rect 338724 3516 338730 3528
rect 339402 3516 339408 3528
rect 338724 3488 339408 3516
rect 338724 3476 338730 3488
rect 339402 3476 339408 3488
rect 339460 3476 339466 3528
rect 340966 3476 340972 3528
rect 341024 3516 341030 3528
rect 341978 3516 341984 3528
rect 341024 3488 341984 3516
rect 341024 3476 341030 3488
rect 341978 3476 341984 3488
rect 342036 3476 342042 3528
rect 348050 3476 348056 3528
rect 348108 3516 348114 3528
rect 349062 3516 349068 3528
rect 348108 3488 349068 3516
rect 348108 3476 348114 3488
rect 349062 3476 349068 3488
rect 349120 3476 349126 3528
rect 349246 3476 349252 3528
rect 349304 3516 349310 3528
rect 350442 3516 350448 3528
rect 349304 3488 350448 3516
rect 349304 3476 349310 3488
rect 350442 3476 350448 3488
rect 350500 3476 350506 3528
rect 355321 3519 355379 3525
rect 355321 3485 355333 3519
rect 355367 3516 355379 3519
rect 404725 3519 404783 3525
rect 404725 3516 404737 3519
rect 355367 3488 404737 3516
rect 355367 3485 355379 3488
rect 355321 3479 355379 3485
rect 404725 3485 404737 3488
rect 404771 3485 404783 3519
rect 404725 3479 404783 3485
rect 404814 3476 404820 3528
rect 404872 3516 404878 3528
rect 405642 3516 405648 3528
rect 404872 3488 405648 3516
rect 404872 3476 404878 3488
rect 405642 3476 405648 3488
rect 405700 3476 405706 3528
rect 406010 3476 406016 3528
rect 406068 3516 406074 3528
rect 407022 3516 407028 3528
rect 406068 3488 407028 3516
rect 406068 3476 406074 3488
rect 407022 3476 407028 3488
rect 407080 3476 407086 3528
rect 407206 3476 407212 3528
rect 407264 3516 407270 3528
rect 409138 3516 409144 3528
rect 407264 3488 409144 3516
rect 407264 3476 407270 3488
rect 409138 3476 409144 3488
rect 409196 3476 409202 3528
rect 409598 3476 409604 3528
rect 409656 3516 409662 3528
rect 410518 3516 410524 3528
rect 409656 3488 410524 3516
rect 409656 3476 409662 3488
rect 410518 3476 410524 3488
rect 410576 3476 410582 3528
rect 411898 3476 411904 3528
rect 411956 3516 411962 3528
rect 412542 3516 412548 3528
rect 411956 3488 412548 3516
rect 411956 3476 411962 3488
rect 412542 3476 412548 3488
rect 412600 3476 412606 3528
rect 413094 3476 413100 3528
rect 413152 3516 413158 3528
rect 413922 3516 413928 3528
rect 413152 3488 413928 3516
rect 413152 3476 413158 3488
rect 413922 3476 413928 3488
rect 413980 3476 413986 3528
rect 414290 3476 414296 3528
rect 414348 3516 414354 3528
rect 415302 3516 415308 3528
rect 414348 3488 415308 3516
rect 414348 3476 414354 3488
rect 415302 3476 415308 3488
rect 415360 3476 415366 3528
rect 416682 3476 416688 3528
rect 416740 3516 416746 3528
rect 417418 3516 417424 3528
rect 416740 3488 417424 3516
rect 416740 3476 416746 3488
rect 417418 3476 417424 3488
rect 417476 3476 417482 3528
rect 418982 3476 418988 3528
rect 419040 3516 419046 3528
rect 419442 3516 419448 3528
rect 419040 3488 419448 3516
rect 419040 3476 419046 3488
rect 419442 3476 419448 3488
rect 419500 3476 419506 3528
rect 419537 3519 419595 3525
rect 419537 3485 419549 3519
rect 419583 3516 419595 3519
rect 461026 3516 461032 3528
rect 419583 3488 461032 3516
rect 419583 3485 419595 3488
rect 419537 3479 419595 3485
rect 461026 3476 461032 3488
rect 461084 3476 461090 3528
rect 471054 3476 471060 3528
rect 471112 3516 471118 3528
rect 471882 3516 471888 3528
rect 471112 3488 471888 3516
rect 471112 3476 471118 3488
rect 471882 3476 471888 3488
rect 471940 3476 471946 3528
rect 478138 3476 478144 3528
rect 478196 3516 478202 3528
rect 479518 3516 479524 3528
rect 478196 3488 479524 3516
rect 478196 3476 478202 3488
rect 479518 3476 479524 3488
rect 479576 3476 479582 3528
rect 480226 3516 480254 3556
rect 481726 3544 481732 3596
rect 481784 3584 481790 3596
rect 482922 3584 482928 3596
rect 481784 3556 482928 3584
rect 481784 3544 481790 3556
rect 482922 3544 482928 3556
rect 482980 3544 482986 3596
rect 485222 3544 485228 3596
rect 485280 3584 485286 3596
rect 485682 3584 485688 3596
rect 485280 3556 485688 3584
rect 485280 3544 485286 3556
rect 485682 3544 485688 3556
rect 485740 3544 485746 3596
rect 486418 3544 486424 3596
rect 486476 3584 486482 3596
rect 487062 3584 487068 3596
rect 486476 3556 487068 3584
rect 486476 3544 486482 3556
rect 487062 3544 487068 3556
rect 487120 3544 487126 3596
rect 487614 3544 487620 3596
rect 487672 3584 487678 3596
rect 489178 3584 489184 3596
rect 487672 3556 489184 3584
rect 487672 3544 487678 3556
rect 489178 3544 489184 3556
rect 489236 3544 489242 3596
rect 489273 3587 489331 3593
rect 489273 3553 489285 3587
rect 489319 3584 489331 3587
rect 504376 3584 504404 3624
rect 510614 3612 510620 3624
rect 510672 3612 510678 3664
rect 519538 3652 519544 3664
rect 514036 3624 519544 3652
rect 489319 3556 504404 3584
rect 489319 3553 489331 3556
rect 489273 3547 489331 3553
rect 505370 3544 505376 3596
rect 505428 3584 505434 3596
rect 514036 3584 514064 3624
rect 519538 3612 519544 3624
rect 519596 3612 519602 3664
rect 535546 3652 535552 3664
rect 528526 3624 535552 3652
rect 505428 3556 514064 3584
rect 505428 3544 505434 3556
rect 518342 3544 518348 3596
rect 518400 3584 518406 3596
rect 528526 3584 528554 3624
rect 535546 3612 535552 3624
rect 535604 3612 535610 3664
rect 554958 3612 554964 3664
rect 555016 3652 555022 3664
rect 558178 3652 558184 3664
rect 555016 3624 558184 3652
rect 555016 3612 555022 3624
rect 558178 3612 558184 3624
rect 558236 3612 558242 3664
rect 566826 3612 566832 3664
rect 566884 3652 566890 3664
rect 570138 3652 570144 3664
rect 566884 3624 570144 3652
rect 566884 3612 566890 3624
rect 570138 3612 570144 3624
rect 570196 3612 570202 3664
rect 518400 3556 528554 3584
rect 518400 3544 518406 3556
rect 533706 3544 533712 3596
rect 533764 3584 533770 3596
rect 546586 3584 546592 3596
rect 533764 3556 546592 3584
rect 533764 3544 533770 3556
rect 546586 3544 546592 3556
rect 546644 3544 546650 3596
rect 546678 3544 546684 3596
rect 546736 3584 546742 3596
rect 548518 3584 548524 3596
rect 546736 3556 548524 3584
rect 546736 3544 546742 3556
rect 548518 3544 548524 3556
rect 548576 3544 548582 3596
rect 551462 3544 551468 3596
rect 551520 3584 551526 3596
rect 556798 3584 556804 3596
rect 551520 3556 556804 3584
rect 551520 3544 551526 3556
rect 556798 3544 556804 3556
rect 556856 3544 556862 3596
rect 559742 3544 559748 3596
rect 559800 3584 559806 3596
rect 565998 3584 566004 3596
rect 559800 3556 566004 3584
rect 559800 3544 559806 3556
rect 565998 3544 566004 3556
rect 566056 3544 566062 3596
rect 570322 3544 570328 3596
rect 570380 3584 570386 3596
rect 572714 3584 572720 3596
rect 570380 3556 572720 3584
rect 570380 3544 570386 3556
rect 572714 3544 572720 3556
rect 572772 3544 572778 3596
rect 501601 3519 501659 3525
rect 501601 3516 501613 3519
rect 480226 3488 501613 3516
rect 501601 3485 501613 3488
rect 501647 3485 501659 3519
rect 501601 3479 501659 3485
rect 501782 3476 501788 3528
rect 501840 3516 501846 3528
rect 502242 3516 502248 3528
rect 501840 3488 502248 3516
rect 501840 3476 501846 3488
rect 502242 3476 502248 3488
rect 502300 3476 502306 3528
rect 502978 3476 502984 3528
rect 503036 3516 503042 3528
rect 503622 3516 503628 3528
rect 503036 3488 503628 3516
rect 503036 3476 503042 3488
rect 503622 3476 503628 3488
rect 503680 3476 503686 3528
rect 507670 3476 507676 3528
rect 507728 3516 507734 3528
rect 528646 3516 528652 3528
rect 507728 3488 528652 3516
rect 507728 3476 507734 3488
rect 528646 3476 528652 3488
rect 528704 3476 528710 3528
rect 529014 3476 529020 3528
rect 529072 3516 529078 3528
rect 529842 3516 529848 3528
rect 529072 3488 529848 3516
rect 529072 3476 529078 3488
rect 529842 3476 529848 3488
rect 529900 3476 529906 3528
rect 532510 3476 532516 3528
rect 532568 3516 532574 3528
rect 533338 3516 533344 3528
rect 532568 3488 533344 3516
rect 532568 3476 532574 3488
rect 533338 3476 533344 3488
rect 533396 3476 533402 3528
rect 534902 3476 534908 3528
rect 534960 3516 534966 3528
rect 535362 3516 535368 3528
rect 534960 3488 535368 3516
rect 534960 3476 534966 3488
rect 535362 3476 535368 3488
rect 535420 3476 535426 3528
rect 536098 3476 536104 3528
rect 536156 3516 536162 3528
rect 536742 3516 536748 3528
rect 536156 3488 536748 3516
rect 536156 3476 536162 3488
rect 536742 3476 536748 3488
rect 536800 3476 536806 3528
rect 537202 3476 537208 3528
rect 537260 3516 537266 3528
rect 538122 3516 538128 3528
rect 537260 3488 538128 3516
rect 537260 3476 537266 3488
rect 538122 3476 538128 3488
rect 538180 3476 538186 3528
rect 538398 3476 538404 3528
rect 538456 3516 538462 3528
rect 539502 3516 539508 3528
rect 538456 3488 539508 3516
rect 538456 3476 538462 3488
rect 539502 3476 539508 3488
rect 539560 3476 539566 3528
rect 541986 3476 541992 3528
rect 542044 3516 542050 3528
rect 542998 3516 543004 3528
rect 542044 3488 543004 3516
rect 542044 3476 542050 3488
rect 542998 3476 543004 3488
rect 543056 3476 543062 3528
rect 543182 3476 543188 3528
rect 543240 3516 543246 3528
rect 544286 3516 544292 3528
rect 543240 3488 544292 3516
rect 543240 3476 543246 3488
rect 544286 3476 544292 3488
rect 544344 3476 544350 3528
rect 544378 3476 544384 3528
rect 544436 3516 544442 3528
rect 545022 3516 545028 3528
rect 544436 3488 545028 3516
rect 544436 3476 544442 3488
rect 545022 3476 545028 3488
rect 545080 3476 545086 3528
rect 545482 3476 545488 3528
rect 545540 3516 545546 3528
rect 547138 3516 547144 3528
rect 545540 3488 547144 3516
rect 545540 3476 545546 3488
rect 547138 3476 547144 3488
rect 547196 3476 547202 3528
rect 550266 3476 550272 3528
rect 550324 3516 550330 3528
rect 551278 3516 551284 3528
rect 550324 3488 551284 3516
rect 550324 3476 550330 3488
rect 551278 3476 551284 3488
rect 551336 3476 551342 3528
rect 553762 3476 553768 3528
rect 553820 3516 553826 3528
rect 554682 3516 554688 3528
rect 553820 3488 554688 3516
rect 553820 3476 553826 3488
rect 554682 3476 554688 3488
rect 554740 3476 554746 3528
rect 560846 3476 560852 3528
rect 560904 3516 560910 3528
rect 561582 3516 561588 3528
rect 560904 3488 561588 3516
rect 560904 3476 560910 3488
rect 561582 3476 561588 3488
rect 561640 3476 561646 3528
rect 562042 3476 562048 3528
rect 562100 3516 562106 3528
rect 562962 3516 562968 3528
rect 562100 3488 562968 3516
rect 562100 3476 562106 3488
rect 562962 3476 562968 3488
rect 563020 3476 563026 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 566458 3516 566464 3528
rect 564492 3488 566464 3516
rect 564492 3476 564498 3488
rect 566458 3476 566464 3488
rect 566516 3476 566522 3528
rect 568022 3476 568028 3528
rect 568080 3516 568086 3528
rect 569218 3516 569224 3528
rect 568080 3488 569224 3516
rect 568080 3476 568086 3488
rect 569218 3476 569224 3488
rect 569276 3476 569282 3528
rect 571518 3476 571524 3528
rect 571576 3516 571582 3528
rect 572622 3516 572628 3528
rect 571576 3488 572628 3516
rect 571576 3476 571582 3488
rect 572622 3476 572628 3488
rect 572680 3476 572686 3528
rect 577406 3476 577412 3528
rect 577464 3516 577470 3528
rect 578234 3516 578240 3528
rect 577464 3488 578240 3516
rect 577464 3476 577470 3488
rect 578234 3476 578240 3488
rect 578292 3476 578298 3528
rect 583021 3519 583079 3525
rect 583021 3485 583033 3519
rect 583067 3516 583079 3519
rect 583386 3516 583392 3528
rect 583067 3488 583392 3516
rect 583067 3485 583079 3488
rect 583021 3479 583079 3485
rect 583386 3476 583392 3488
rect 583444 3476 583450 3528
rect 238018 3448 238024 3460
rect 186188 3420 222516 3448
rect 222672 3420 238024 3448
rect 186188 3408 186194 3420
rect 23014 3340 23020 3392
rect 23072 3380 23078 3392
rect 38289 3383 38347 3389
rect 38289 3380 38301 3383
rect 23072 3352 38301 3380
rect 23072 3340 23078 3352
rect 38289 3349 38301 3352
rect 38335 3349 38347 3383
rect 40773 3383 40831 3389
rect 40773 3380 40785 3383
rect 38289 3343 38347 3349
rect 39500 3352 40785 3380
rect 6454 3272 6460 3324
rect 6512 3312 6518 3324
rect 7558 3312 7564 3324
rect 6512 3284 7564 3312
rect 6512 3272 6518 3284
rect 7558 3272 7564 3284
rect 7616 3272 7622 3324
rect 24210 3272 24216 3324
rect 24268 3312 24274 3324
rect 24268 3284 26234 3312
rect 24268 3272 24274 3284
rect 26206 3244 26234 3284
rect 31294 3272 31300 3324
rect 31352 3312 31358 3324
rect 39500 3312 39528 3352
rect 40773 3349 40785 3352
rect 40819 3349 40831 3383
rect 40773 3343 40831 3349
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 58618 3380 58624 3392
rect 41932 3352 58624 3380
rect 41932 3340 41938 3352
rect 58618 3340 58624 3352
rect 58676 3340 58682 3392
rect 74994 3340 75000 3392
rect 75052 3380 75058 3392
rect 196618 3380 196624 3392
rect 75052 3352 196624 3380
rect 75052 3340 75058 3352
rect 196618 3340 196624 3352
rect 196676 3340 196682 3392
rect 219250 3340 219256 3392
rect 219308 3380 219314 3392
rect 219308 3352 219434 3380
rect 219308 3340 219314 3352
rect 31352 3284 39528 3312
rect 31352 3272 31358 3284
rect 39574 3272 39580 3324
rect 39632 3312 39638 3324
rect 43438 3312 43444 3324
rect 39632 3284 43444 3312
rect 39632 3272 39638 3284
rect 43438 3272 43444 3284
rect 43496 3272 43502 3324
rect 45462 3272 45468 3324
rect 45520 3312 45526 3324
rect 61378 3312 61384 3324
rect 45520 3284 61384 3312
rect 45520 3272 45526 3284
rect 61378 3272 61384 3284
rect 61436 3272 61442 3324
rect 80882 3272 80888 3324
rect 80940 3312 80946 3324
rect 81342 3312 81348 3324
rect 80940 3284 81348 3312
rect 80940 3272 80946 3284
rect 81342 3272 81348 3284
rect 81400 3272 81406 3324
rect 84470 3272 84476 3324
rect 84528 3312 84534 3324
rect 85482 3312 85488 3324
rect 84528 3284 85488 3312
rect 84528 3272 84534 3284
rect 85482 3272 85488 3284
rect 85540 3272 85546 3324
rect 85577 3315 85635 3321
rect 85577 3281 85589 3315
rect 85623 3312 85635 3315
rect 87598 3312 87604 3324
rect 85623 3284 87604 3312
rect 85623 3281 85635 3284
rect 85577 3275 85635 3281
rect 87598 3272 87604 3284
rect 87656 3272 87662 3324
rect 87966 3272 87972 3324
rect 88024 3312 88030 3324
rect 88978 3312 88984 3324
rect 88024 3284 88984 3312
rect 88024 3272 88030 3284
rect 88978 3272 88984 3284
rect 89036 3272 89042 3324
rect 199378 3312 199384 3324
rect 89088 3284 199384 3312
rect 35158 3244 35164 3256
rect 26206 3216 35164 3244
rect 35158 3204 35164 3216
rect 35216 3204 35222 3256
rect 38289 3247 38347 3253
rect 38289 3213 38301 3247
rect 38335 3244 38347 3247
rect 40678 3244 40684 3256
rect 38335 3216 40684 3244
rect 38335 3213 38347 3216
rect 38289 3207 38347 3213
rect 40678 3204 40684 3216
rect 40736 3204 40742 3256
rect 82078 3204 82084 3256
rect 82136 3244 82142 3256
rect 89088 3244 89116 3284
rect 199378 3272 199384 3284
rect 199436 3272 199442 3324
rect 82136 3216 89116 3244
rect 82136 3204 82142 3216
rect 91554 3204 91560 3256
rect 91612 3244 91618 3256
rect 93118 3244 93124 3256
rect 91612 3216 93124 3244
rect 91612 3204 91618 3216
rect 93118 3204 93124 3216
rect 93176 3204 93182 3256
rect 200758 3244 200764 3256
rect 93228 3216 200764 3244
rect 15930 3136 15936 3188
rect 15988 3176 15994 3188
rect 17218 3176 17224 3188
rect 15988 3148 17224 3176
rect 15988 3136 15994 3148
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 50154 3136 50160 3188
rect 50212 3176 50218 3188
rect 86218 3176 86224 3188
rect 50212 3148 86224 3176
rect 50212 3136 50218 3148
rect 86218 3136 86224 3148
rect 86276 3136 86282 3188
rect 57238 3068 57244 3120
rect 57296 3108 57302 3120
rect 85577 3111 85635 3117
rect 85577 3108 85589 3111
rect 57296 3080 85589 3108
rect 57296 3068 57302 3080
rect 85577 3077 85589 3080
rect 85623 3077 85635 3111
rect 85577 3071 85635 3077
rect 85666 3068 85672 3120
rect 85724 3108 85730 3120
rect 93228 3108 93256 3216
rect 200758 3204 200764 3216
rect 200816 3204 200822 3256
rect 219406 3244 219434 3352
rect 222488 3312 222516 3420
rect 238018 3408 238024 3420
rect 238076 3408 238082 3460
rect 238110 3408 238116 3460
rect 238168 3448 238174 3460
rect 326709 3451 326767 3457
rect 326709 3448 326721 3451
rect 238168 3420 326721 3448
rect 238168 3408 238174 3420
rect 326709 3417 326721 3420
rect 326755 3417 326767 3451
rect 326709 3411 326767 3417
rect 326798 3408 326804 3460
rect 326856 3448 326862 3460
rect 329098 3448 329104 3460
rect 326856 3420 329104 3448
rect 326856 3408 326862 3420
rect 329098 3408 329104 3420
rect 329156 3408 329162 3460
rect 331582 3408 331588 3460
rect 331640 3448 331646 3460
rect 332502 3448 332508 3460
rect 331640 3420 332508 3448
rect 331640 3408 331646 3420
rect 332502 3408 332508 3420
rect 332560 3408 332566 3460
rect 337470 3408 337476 3460
rect 337528 3448 337534 3460
rect 405826 3448 405832 3460
rect 337528 3420 405832 3448
rect 337528 3408 337534 3420
rect 405826 3408 405832 3420
rect 405884 3408 405890 3460
rect 408402 3408 408408 3460
rect 408460 3448 408466 3460
rect 451277 3451 451335 3457
rect 451277 3448 451289 3451
rect 408460 3420 451289 3448
rect 408460 3408 408466 3420
rect 451277 3417 451289 3420
rect 451323 3417 451335 3451
rect 456058 3448 456064 3460
rect 451277 3411 451335 3417
rect 451384 3420 456064 3448
rect 231118 3380 231124 3392
rect 224926 3352 231124 3380
rect 224926 3312 224954 3352
rect 231118 3340 231124 3352
rect 231176 3340 231182 3392
rect 237374 3380 237380 3392
rect 231228 3352 237380 3380
rect 222488 3284 224954 3312
rect 226334 3272 226340 3324
rect 226392 3312 226398 3324
rect 227622 3312 227628 3324
rect 226392 3284 227628 3312
rect 226392 3272 226398 3284
rect 227622 3272 227628 3284
rect 227680 3272 227686 3324
rect 219406 3216 224954 3244
rect 203518 3176 203524 3188
rect 93826 3148 203524 3176
rect 85724 3080 93256 3108
rect 85724 3068 85730 3080
rect 93302 3068 93308 3120
rect 93360 3108 93366 3120
rect 93826 3108 93854 3148
rect 203518 3136 203524 3148
rect 203576 3136 203582 3188
rect 224926 3176 224954 3216
rect 231228 3176 231256 3352
rect 237374 3340 237380 3352
rect 237432 3340 237438 3392
rect 240502 3340 240508 3392
rect 240560 3380 240566 3392
rect 267826 3380 267832 3392
rect 240560 3352 267832 3380
rect 240560 3340 240566 3352
rect 267826 3340 267832 3352
rect 267884 3340 267890 3392
rect 270034 3340 270040 3392
rect 270092 3380 270098 3392
rect 298373 3383 298431 3389
rect 298373 3380 298385 3383
rect 270092 3352 298385 3380
rect 270092 3340 270098 3352
rect 298373 3349 298385 3352
rect 298419 3349 298431 3383
rect 298373 3343 298431 3349
rect 298462 3340 298468 3392
rect 298520 3380 298526 3392
rect 299382 3380 299388 3392
rect 298520 3352 299388 3380
rect 298520 3340 298526 3352
rect 299382 3340 299388 3352
rect 299440 3340 299446 3392
rect 305546 3340 305552 3392
rect 305604 3380 305610 3392
rect 306282 3380 306288 3392
rect 305604 3352 306288 3380
rect 305604 3340 305610 3352
rect 306282 3340 306288 3352
rect 306340 3340 306346 3392
rect 312630 3340 312636 3392
rect 312688 3380 312694 3392
rect 313182 3380 313188 3392
rect 312688 3352 313188 3380
rect 312688 3340 312694 3352
rect 313182 3340 313188 3352
rect 313240 3340 313246 3392
rect 323302 3340 323308 3392
rect 323360 3380 323366 3392
rect 325053 3383 325111 3389
rect 325053 3380 325065 3383
rect 323360 3352 325065 3380
rect 323360 3340 323366 3352
rect 325053 3349 325065 3352
rect 325099 3349 325111 3383
rect 325053 3343 325111 3349
rect 329190 3340 329196 3392
rect 329248 3380 329254 3392
rect 331858 3380 331864 3392
rect 329248 3352 331864 3380
rect 329248 3340 329254 3352
rect 331858 3340 331864 3352
rect 331916 3340 331922 3392
rect 350442 3340 350448 3392
rect 350500 3380 350506 3392
rect 352558 3380 352564 3392
rect 350500 3352 352564 3380
rect 350500 3340 350506 3352
rect 352558 3340 352564 3352
rect 352616 3340 352622 3392
rect 354677 3383 354735 3389
rect 354677 3349 354689 3383
rect 354723 3380 354735 3383
rect 358814 3380 358820 3392
rect 354723 3352 358820 3380
rect 354723 3349 354735 3352
rect 354677 3343 354735 3349
rect 358814 3340 358820 3352
rect 358872 3340 358878 3392
rect 363506 3340 363512 3392
rect 363564 3380 363570 3392
rect 364242 3380 364248 3392
rect 363564 3352 364248 3380
rect 363564 3340 363570 3352
rect 364242 3340 364248 3352
rect 364300 3340 364306 3392
rect 364610 3340 364616 3392
rect 364668 3380 364674 3392
rect 366358 3380 366364 3392
rect 364668 3352 366364 3380
rect 364668 3340 364674 3352
rect 366358 3340 366364 3352
rect 366416 3340 366422 3392
rect 367002 3340 367008 3392
rect 367060 3380 367066 3392
rect 367738 3380 367744 3392
rect 367060 3352 367744 3380
rect 367060 3340 367066 3352
rect 367738 3340 367744 3352
rect 367796 3340 367802 3392
rect 371694 3340 371700 3392
rect 371752 3380 371758 3392
rect 373258 3380 373264 3392
rect 371752 3352 373264 3380
rect 371752 3340 371758 3352
rect 373258 3340 373264 3352
rect 373316 3340 373322 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 376478 3340 376484 3392
rect 376536 3380 376542 3392
rect 377398 3380 377404 3392
rect 376536 3352 377404 3380
rect 376536 3340 376542 3352
rect 377398 3340 377404 3352
rect 377456 3340 377462 3392
rect 378870 3340 378876 3392
rect 378928 3380 378934 3392
rect 379422 3380 379428 3392
rect 378928 3352 379428 3380
rect 378928 3340 378934 3352
rect 379422 3340 379428 3352
rect 379480 3340 379486 3392
rect 381170 3340 381176 3392
rect 381228 3380 381234 3392
rect 382918 3380 382924 3392
rect 381228 3352 382924 3380
rect 381228 3340 381234 3352
rect 382918 3340 382924 3352
rect 382976 3340 382982 3392
rect 383013 3383 383071 3389
rect 383013 3349 383025 3383
rect 383059 3380 383071 3383
rect 423677 3383 423735 3389
rect 423677 3380 423689 3383
rect 383059 3352 423689 3380
rect 383059 3349 383071 3352
rect 383013 3343 383071 3349
rect 423677 3349 423689 3352
rect 423723 3349 423735 3383
rect 423677 3343 423735 3349
rect 423766 3340 423772 3392
rect 423824 3380 423830 3392
rect 425790 3380 425796 3392
rect 423824 3352 425796 3380
rect 423824 3340 423830 3352
rect 425790 3340 425796 3352
rect 425848 3340 425854 3392
rect 427262 3340 427268 3392
rect 427320 3380 427326 3392
rect 428458 3380 428464 3392
rect 427320 3352 428464 3380
rect 427320 3340 427326 3352
rect 428458 3340 428464 3352
rect 428516 3340 428522 3392
rect 429654 3340 429660 3392
rect 429712 3380 429718 3392
rect 430482 3380 430488 3392
rect 429712 3352 430488 3380
rect 429712 3340 429718 3352
rect 430482 3340 430488 3352
rect 430540 3340 430546 3392
rect 430850 3340 430856 3392
rect 430908 3380 430914 3392
rect 431862 3380 431868 3392
rect 430908 3352 431868 3380
rect 430908 3340 430914 3352
rect 431862 3340 431868 3352
rect 431920 3340 431926 3392
rect 432046 3340 432052 3392
rect 432104 3380 432110 3392
rect 433242 3380 433248 3392
rect 432104 3352 433248 3380
rect 432104 3340 432110 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 436646 3380 436652 3392
rect 434272 3352 436652 3380
rect 233418 3272 233424 3324
rect 233476 3312 233482 3324
rect 258166 3312 258172 3324
rect 233476 3284 258172 3312
rect 233476 3272 233482 3284
rect 258166 3272 258172 3284
rect 258224 3272 258230 3324
rect 258258 3272 258264 3324
rect 258316 3312 258322 3324
rect 260098 3312 260104 3324
rect 258316 3284 260104 3312
rect 258316 3272 258322 3284
rect 260098 3272 260104 3284
rect 260156 3272 260162 3324
rect 277118 3272 277124 3324
rect 277176 3312 277182 3324
rect 307018 3312 307024 3324
rect 277176 3284 307024 3312
rect 277176 3272 277182 3284
rect 307018 3272 307024 3284
rect 307076 3272 307082 3324
rect 309042 3272 309048 3324
rect 309100 3312 309106 3324
rect 385034 3312 385040 3324
rect 309100 3284 385040 3312
rect 309100 3272 309106 3284
rect 385034 3272 385040 3284
rect 385092 3272 385098 3324
rect 388254 3272 388260 3324
rect 388312 3312 388318 3324
rect 389910 3312 389916 3324
rect 388312 3284 389916 3312
rect 388312 3272 388318 3284
rect 389910 3272 389916 3284
rect 389968 3272 389974 3324
rect 390646 3272 390652 3324
rect 390704 3312 390710 3324
rect 391750 3312 391756 3324
rect 390704 3284 391756 3312
rect 390704 3272 390710 3284
rect 391750 3272 391756 3284
rect 391808 3272 391814 3324
rect 391842 3272 391848 3324
rect 391900 3312 391906 3324
rect 392578 3312 392584 3324
rect 391900 3284 392584 3312
rect 391900 3272 391906 3284
rect 392578 3272 392584 3284
rect 392636 3272 392642 3324
rect 392673 3315 392731 3321
rect 392673 3281 392685 3315
rect 392719 3312 392731 3315
rect 434272 3312 434300 3352
rect 436646 3340 436652 3352
rect 436704 3340 436710 3392
rect 436738 3340 436744 3392
rect 436796 3380 436802 3392
rect 437382 3380 437388 3392
rect 436796 3352 437388 3380
rect 436796 3340 436802 3352
rect 437382 3340 437388 3352
rect 437440 3340 437446 3392
rect 439130 3340 439136 3392
rect 439188 3380 439194 3392
rect 440142 3380 440148 3392
rect 439188 3352 440148 3380
rect 439188 3340 439194 3352
rect 440142 3340 440148 3352
rect 440200 3340 440206 3392
rect 440237 3383 440295 3389
rect 440237 3349 440249 3383
rect 440283 3380 440295 3383
rect 451384 3380 451412 3420
rect 456058 3408 456064 3420
rect 456116 3408 456122 3460
rect 460382 3408 460388 3460
rect 460440 3448 460446 3460
rect 462958 3448 462964 3460
rect 460440 3420 462964 3448
rect 460440 3408 460446 3420
rect 462958 3408 462964 3420
rect 463016 3408 463022 3460
rect 463970 3408 463976 3460
rect 464028 3448 464034 3460
rect 464028 3420 492260 3448
rect 464028 3408 464034 3420
rect 440283 3352 451412 3380
rect 440283 3349 440295 3352
rect 440237 3343 440295 3349
rect 452102 3340 452108 3392
rect 452160 3380 452166 3392
rect 453298 3380 453304 3392
rect 452160 3352 453304 3380
rect 452160 3340 452166 3352
rect 453298 3340 453304 3352
rect 453356 3340 453362 3392
rect 456978 3380 456984 3392
rect 453408 3352 456984 3380
rect 392719 3284 434300 3312
rect 392719 3281 392731 3284
rect 392673 3275 392731 3281
rect 434438 3272 434444 3324
rect 434496 3312 434502 3324
rect 435358 3312 435364 3324
rect 434496 3284 435364 3312
rect 434496 3272 434502 3284
rect 435358 3272 435364 3284
rect 435416 3272 435422 3324
rect 435453 3315 435511 3321
rect 435453 3281 435465 3315
rect 435499 3312 435511 3315
rect 437753 3315 437811 3321
rect 437753 3312 437765 3315
rect 435499 3284 437765 3312
rect 435499 3281 435511 3284
rect 435453 3275 435511 3281
rect 437753 3281 437765 3284
rect 437799 3281 437811 3315
rect 437753 3275 437811 3281
rect 437934 3272 437940 3324
rect 437992 3312 437998 3324
rect 440878 3312 440884 3324
rect 437992 3284 440884 3312
rect 437992 3272 437998 3284
rect 440878 3272 440884 3284
rect 440936 3272 440942 3324
rect 441522 3272 441528 3324
rect 441580 3312 441586 3324
rect 446398 3312 446404 3324
rect 441580 3284 446404 3312
rect 441580 3272 441586 3284
rect 446398 3272 446404 3284
rect 446456 3272 446462 3324
rect 447410 3272 447416 3324
rect 447468 3312 447474 3324
rect 450633 3315 450691 3321
rect 450633 3312 450645 3315
rect 447468 3284 450645 3312
rect 447468 3272 447474 3284
rect 450633 3281 450645 3284
rect 450679 3281 450691 3315
rect 450633 3275 450691 3281
rect 451277 3315 451335 3321
rect 451277 3281 451289 3315
rect 451323 3312 451335 3315
rect 453408 3312 453436 3352
rect 456978 3340 456984 3352
rect 457036 3340 457042 3392
rect 461578 3340 461584 3392
rect 461636 3380 461642 3392
rect 471517 3383 471575 3389
rect 471517 3380 471529 3383
rect 461636 3352 471529 3380
rect 461636 3340 461642 3352
rect 471517 3349 471529 3352
rect 471563 3349 471575 3383
rect 472710 3380 472716 3392
rect 471517 3343 471575 3349
rect 471624 3352 472716 3380
rect 451323 3284 453436 3312
rect 451323 3281 451335 3284
rect 451277 3275 451335 3281
rect 455690 3272 455696 3324
rect 455748 3312 455754 3324
rect 471624 3312 471652 3352
rect 472710 3340 472716 3352
rect 472768 3340 472774 3392
rect 480530 3340 480536 3392
rect 480588 3380 480594 3392
rect 482278 3380 482284 3392
rect 480588 3352 482284 3380
rect 480588 3340 480594 3352
rect 482278 3340 482284 3352
rect 482336 3340 482342 3392
rect 488810 3340 488816 3392
rect 488868 3380 488874 3392
rect 489822 3380 489828 3392
rect 488868 3352 489828 3380
rect 488868 3340 488874 3352
rect 489822 3340 489828 3352
rect 489880 3340 489886 3392
rect 492232 3380 492260 3420
rect 492306 3408 492312 3460
rect 492364 3448 492370 3460
rect 493318 3448 493324 3460
rect 492364 3420 493324 3448
rect 492364 3408 492370 3420
rect 493318 3408 493324 3420
rect 493376 3408 493382 3460
rect 494698 3408 494704 3460
rect 494756 3448 494762 3460
rect 495342 3448 495348 3460
rect 494756 3420 495348 3448
rect 494756 3408 494762 3420
rect 495342 3408 495348 3420
rect 495400 3408 495406 3460
rect 495894 3408 495900 3460
rect 495952 3448 495958 3460
rect 496722 3448 496728 3460
rect 495952 3420 496728 3448
rect 495952 3408 495958 3420
rect 496722 3408 496728 3420
rect 496780 3408 496786 3460
rect 499390 3408 499396 3460
rect 499448 3448 499454 3460
rect 499448 3420 509234 3448
rect 499448 3408 499454 3420
rect 496998 3380 497004 3392
rect 492232 3352 497004 3380
rect 496998 3340 497004 3352
rect 497056 3340 497062 3392
rect 509206 3380 509234 3420
rect 511258 3408 511264 3460
rect 511316 3448 511322 3460
rect 511902 3448 511908 3460
rect 511316 3420 511908 3448
rect 511316 3408 511322 3420
rect 511902 3408 511908 3420
rect 511960 3408 511966 3460
rect 512454 3408 512460 3460
rect 512512 3448 512518 3460
rect 513282 3448 513288 3460
rect 512512 3420 513288 3448
rect 512512 3408 512518 3420
rect 513282 3408 513288 3420
rect 513340 3408 513346 3460
rect 513558 3408 513564 3460
rect 513616 3448 513622 3460
rect 514662 3448 514668 3460
rect 513616 3420 514668 3448
rect 513616 3408 513622 3420
rect 514662 3408 514668 3420
rect 514720 3408 514726 3460
rect 514754 3408 514760 3460
rect 514812 3448 514818 3460
rect 515858 3448 515864 3460
rect 514812 3420 515864 3448
rect 514812 3408 514818 3420
rect 515858 3408 515864 3420
rect 515916 3408 515922 3460
rect 519538 3408 519544 3460
rect 519596 3448 519602 3460
rect 520182 3448 520188 3460
rect 519596 3420 520188 3448
rect 519596 3408 519602 3420
rect 520182 3408 520188 3420
rect 520240 3408 520246 3460
rect 520734 3408 520740 3460
rect 520792 3448 520798 3460
rect 521562 3448 521568 3460
rect 520792 3420 521568 3448
rect 520792 3408 520798 3420
rect 521562 3408 521568 3420
rect 521620 3408 521626 3460
rect 521838 3408 521844 3460
rect 521896 3448 521902 3460
rect 522942 3448 522948 3460
rect 521896 3420 522948 3448
rect 521896 3408 521902 3420
rect 522942 3408 522948 3420
rect 523000 3408 523006 3460
rect 524230 3408 524236 3460
rect 524288 3448 524294 3460
rect 525150 3448 525156 3460
rect 524288 3420 525156 3448
rect 524288 3408 524294 3420
rect 525150 3408 525156 3420
rect 525208 3408 525214 3460
rect 526622 3408 526628 3460
rect 526680 3448 526686 3460
rect 527082 3448 527088 3460
rect 526680 3420 527088 3448
rect 526680 3408 526686 3420
rect 527082 3408 527088 3420
rect 527140 3408 527146 3460
rect 527818 3408 527824 3460
rect 527876 3448 527882 3460
rect 542354 3448 542360 3460
rect 527876 3420 542360 3448
rect 527876 3408 527882 3420
rect 542354 3408 542360 3420
rect 542412 3408 542418 3460
rect 552658 3408 552664 3460
rect 552716 3448 552722 3460
rect 560386 3448 560392 3460
rect 552716 3420 560392 3448
rect 552716 3408 552722 3420
rect 560386 3408 560392 3420
rect 560444 3408 560450 3460
rect 576302 3408 576308 3460
rect 576360 3448 576366 3460
rect 576762 3448 576768 3460
rect 576360 3420 576768 3448
rect 576360 3408 576366 3420
rect 576762 3408 576768 3420
rect 576820 3408 576826 3460
rect 521930 3380 521936 3392
rect 509206 3352 521936 3380
rect 521930 3340 521936 3352
rect 521988 3340 521994 3392
rect 523034 3340 523040 3392
rect 523092 3380 523098 3392
rect 525058 3380 525064 3392
rect 523092 3352 525064 3380
rect 523092 3340 523098 3352
rect 525058 3340 525064 3352
rect 525116 3340 525122 3392
rect 531314 3340 531320 3392
rect 531372 3380 531378 3392
rect 533430 3380 533436 3392
rect 531372 3352 533436 3380
rect 531372 3340 531378 3352
rect 533430 3340 533436 3352
rect 533488 3340 533494 3392
rect 455748 3284 471652 3312
rect 455748 3272 455754 3284
rect 472250 3272 472256 3324
rect 472308 3312 472314 3324
rect 478046 3312 478052 3324
rect 472308 3284 478052 3312
rect 472308 3272 472314 3284
rect 478046 3272 478052 3284
rect 478104 3272 478110 3324
rect 482830 3272 482836 3324
rect 482888 3312 482894 3324
rect 489273 3315 489331 3321
rect 489273 3312 489285 3315
rect 482888 3284 489285 3312
rect 482888 3272 482894 3284
rect 489273 3281 489285 3284
rect 489319 3281 489331 3315
rect 489273 3275 489331 3281
rect 510062 3272 510068 3324
rect 510120 3312 510126 3324
rect 518158 3312 518164 3324
rect 510120 3284 518164 3312
rect 510120 3272 510126 3284
rect 518158 3272 518164 3284
rect 518216 3272 518222 3324
rect 235810 3204 235816 3256
rect 235868 3244 235874 3256
rect 238941 3247 238999 3253
rect 235868 3216 238754 3244
rect 235868 3204 235874 3216
rect 224926 3148 231256 3176
rect 232222 3136 232228 3188
rect 232280 3176 232286 3188
rect 233142 3176 233148 3188
rect 232280 3148 233148 3176
rect 232280 3136 232286 3148
rect 233142 3136 233148 3148
rect 233200 3136 233206 3188
rect 238726 3176 238754 3216
rect 238941 3213 238953 3247
rect 238987 3244 238999 3247
rect 245010 3244 245016 3256
rect 238987 3216 245016 3244
rect 238987 3213 238999 3216
rect 238941 3207 238999 3213
rect 245010 3204 245016 3216
rect 245068 3204 245074 3256
rect 255866 3204 255872 3256
rect 255924 3244 255930 3256
rect 323578 3244 323584 3256
rect 255924 3216 323584 3244
rect 255924 3204 255930 3216
rect 323578 3204 323584 3216
rect 323636 3204 323642 3256
rect 330386 3204 330392 3256
rect 330444 3244 330450 3256
rect 396721 3247 396779 3253
rect 396721 3244 396733 3247
rect 330444 3216 396733 3244
rect 330444 3204 330450 3216
rect 396721 3213 396733 3216
rect 396767 3213 396779 3247
rect 396721 3207 396779 3213
rect 398926 3204 398932 3256
rect 398984 3244 398990 3256
rect 400858 3244 400864 3256
rect 398984 3216 400864 3244
rect 398984 3204 398990 3216
rect 400858 3204 400864 3216
rect 400916 3204 400922 3256
rect 403618 3204 403624 3256
rect 403676 3244 403682 3256
rect 452654 3244 452660 3256
rect 403676 3216 452660 3244
rect 403676 3204 403682 3216
rect 452654 3204 452660 3216
rect 452712 3204 452718 3256
rect 453298 3204 453304 3256
rect 453356 3244 453362 3256
rect 460290 3244 460296 3256
rect 453356 3216 460296 3244
rect 453356 3204 453362 3216
rect 460290 3204 460296 3216
rect 460348 3204 460354 3256
rect 506474 3204 506480 3256
rect 506532 3244 506538 3256
rect 507762 3244 507768 3256
rect 506532 3216 507768 3244
rect 506532 3204 506538 3216
rect 507762 3204 507768 3216
rect 507820 3204 507826 3256
rect 242158 3176 242164 3188
rect 238726 3148 242164 3176
rect 242158 3136 242164 3148
rect 242216 3136 242222 3188
rect 249978 3136 249984 3188
rect 250036 3176 250042 3188
rect 258074 3176 258080 3188
rect 250036 3148 258080 3176
rect 250036 3136 250042 3148
rect 258074 3136 258080 3148
rect 258132 3136 258138 3188
rect 262950 3136 262956 3188
rect 263008 3176 263014 3188
rect 320818 3176 320824 3188
rect 263008 3148 320824 3176
rect 263008 3136 263014 3148
rect 320818 3136 320824 3148
rect 320876 3136 320882 3188
rect 325602 3136 325608 3188
rect 325660 3176 325666 3188
rect 340138 3176 340144 3188
rect 325660 3148 340144 3176
rect 325660 3136 325666 3148
rect 340138 3136 340144 3148
rect 340196 3136 340202 3188
rect 344554 3136 344560 3188
rect 344612 3176 344618 3188
rect 407758 3176 407764 3188
rect 344612 3148 407764 3176
rect 344612 3136 344618 3148
rect 407758 3136 407764 3148
rect 407816 3136 407822 3188
rect 410794 3136 410800 3188
rect 410852 3176 410858 3188
rect 454770 3176 454776 3188
rect 410852 3148 454776 3176
rect 410852 3136 410858 3148
rect 454770 3136 454776 3148
rect 454828 3136 454834 3188
rect 465166 3136 465172 3188
rect 465224 3176 465230 3188
rect 466362 3176 466368 3188
rect 465224 3148 466368 3176
rect 465224 3136 465230 3148
rect 466362 3136 466368 3148
rect 466420 3136 466426 3188
rect 469858 3136 469864 3188
rect 469916 3176 469922 3188
rect 471238 3176 471244 3188
rect 469916 3148 471244 3176
rect 469916 3136 469922 3148
rect 471238 3136 471244 3148
rect 471296 3136 471302 3188
rect 530118 3136 530124 3188
rect 530176 3176 530182 3188
rect 531222 3176 531228 3188
rect 530176 3148 531228 3176
rect 530176 3136 530182 3148
rect 531222 3136 531228 3148
rect 531280 3136 531286 3188
rect 569126 3136 569132 3188
rect 569184 3176 569190 3188
rect 572898 3176 572904 3188
rect 569184 3148 572904 3176
rect 569184 3136 569190 3148
rect 572898 3136 572904 3148
rect 572956 3136 572962 3188
rect 93360 3080 93854 3108
rect 93360 3068 93366 3080
rect 98638 3068 98644 3120
rect 98696 3108 98702 3120
rect 99282 3108 99288 3120
rect 98696 3080 99288 3108
rect 98696 3068 98702 3080
rect 99282 3068 99288 3080
rect 99340 3068 99346 3120
rect 102226 3068 102232 3120
rect 102284 3108 102290 3120
rect 105538 3108 105544 3120
rect 102284 3080 105544 3108
rect 102284 3068 102290 3080
rect 105538 3068 105544 3080
rect 105596 3068 105602 3120
rect 105722 3068 105728 3120
rect 105780 3108 105786 3120
rect 106182 3108 106188 3120
rect 105780 3080 106188 3108
rect 105780 3068 105786 3080
rect 106182 3068 106188 3080
rect 106240 3068 106246 3120
rect 110506 3068 110512 3120
rect 110564 3108 110570 3120
rect 111702 3108 111708 3120
rect 110564 3080 111708 3108
rect 110564 3068 110570 3080
rect 111702 3068 111708 3080
rect 111760 3068 111766 3120
rect 112806 3068 112812 3120
rect 112864 3108 112870 3120
rect 115106 3108 115112 3120
rect 112864 3080 115112 3108
rect 112864 3068 112870 3080
rect 115106 3068 115112 3080
rect 115164 3068 115170 3120
rect 116394 3068 116400 3120
rect 116452 3108 116458 3120
rect 117222 3108 117228 3120
rect 116452 3080 117228 3108
rect 116452 3068 116458 3080
rect 117222 3068 117228 3080
rect 117280 3068 117286 3120
rect 117590 3068 117596 3120
rect 117648 3108 117654 3120
rect 118602 3108 118608 3120
rect 117648 3080 118608 3108
rect 117648 3068 117654 3080
rect 118602 3068 118608 3080
rect 118660 3068 118666 3120
rect 118697 3111 118755 3117
rect 118697 3077 118709 3111
rect 118743 3108 118755 3111
rect 214558 3108 214564 3120
rect 118743 3080 214564 3108
rect 118743 3077 118755 3080
rect 118697 3071 118755 3077
rect 214558 3068 214564 3080
rect 214616 3068 214622 3120
rect 244090 3068 244096 3120
rect 244148 3108 244154 3120
rect 266998 3108 267004 3120
rect 244148 3080 267004 3108
rect 244148 3068 244154 3080
rect 266998 3068 267004 3080
rect 267056 3068 267062 3120
rect 268838 3068 268844 3120
rect 268896 3108 268902 3120
rect 280798 3108 280804 3120
rect 268896 3080 280804 3108
rect 268896 3068 268902 3080
rect 280798 3068 280804 3080
rect 280856 3068 280862 3120
rect 284294 3068 284300 3120
rect 284352 3108 284358 3120
rect 298281 3111 298339 3117
rect 298281 3108 298293 3111
rect 284352 3080 298293 3108
rect 284352 3068 284358 3080
rect 298281 3077 298293 3080
rect 298327 3077 298339 3111
rect 298281 3071 298339 3077
rect 298373 3111 298431 3117
rect 298373 3077 298385 3111
rect 298419 3108 298431 3111
rect 300118 3108 300124 3120
rect 298419 3080 300124 3108
rect 298419 3077 298431 3080
rect 298373 3071 298431 3077
rect 300118 3068 300124 3080
rect 300176 3068 300182 3120
rect 302237 3111 302295 3117
rect 302237 3077 302249 3111
rect 302283 3108 302295 3111
rect 302283 3080 302464 3108
rect 302283 3077 302295 3080
rect 302237 3071 302295 3077
rect 71498 3000 71504 3052
rect 71556 3040 71562 3052
rect 106918 3040 106924 3052
rect 71556 3012 106924 3040
rect 71556 3000 71562 3012
rect 106918 3000 106924 3012
rect 106976 3000 106982 3052
rect 109310 3000 109316 3052
rect 109368 3040 109374 3052
rect 112438 3040 112444 3052
rect 109368 3012 112444 3040
rect 109368 3000 109374 3012
rect 112438 3000 112444 3012
rect 112496 3000 112502 3052
rect 114002 3000 114008 3052
rect 114060 3040 114066 3052
rect 221458 3040 221464 3052
rect 114060 3012 221464 3040
rect 114060 3000 114066 3012
rect 221458 3000 221464 3012
rect 221516 3000 221522 3052
rect 251174 3000 251180 3052
rect 251232 3040 251238 3052
rect 258718 3040 258724 3052
rect 251232 3012 258724 3040
rect 251232 3000 251238 3012
rect 258718 3000 258724 3012
rect 258776 3000 258782 3052
rect 276014 3000 276020 3052
rect 276072 3040 276078 3052
rect 284938 3040 284944 3052
rect 276072 3012 284944 3040
rect 276072 3000 276078 3012
rect 284938 3000 284944 3012
rect 284996 3000 285002 3052
rect 286594 3000 286600 3052
rect 286652 3040 286658 3052
rect 289078 3040 289084 3052
rect 286652 3012 289084 3040
rect 286652 3000 286658 3012
rect 289078 3000 289084 3012
rect 289136 3000 289142 3052
rect 290182 3000 290188 3052
rect 290240 3040 290246 3052
rect 292482 3040 292488 3052
rect 290240 3012 292488 3040
rect 290240 3000 290246 3012
rect 292482 3000 292488 3012
rect 292540 3000 292546 3052
rect 293678 3000 293684 3052
rect 293736 3040 293742 3052
rect 302436 3040 302464 3080
rect 311434 3068 311440 3120
rect 311492 3108 311498 3120
rect 326709 3111 326767 3117
rect 311492 3080 325694 3108
rect 311492 3068 311498 3080
rect 314010 3040 314016 3052
rect 293736 3012 302372 3040
rect 302436 3012 314016 3040
rect 293736 3000 293742 3012
rect 64322 2932 64328 2984
rect 64380 2972 64386 2984
rect 64380 2944 87276 2972
rect 64380 2932 64386 2944
rect 46658 2864 46664 2916
rect 46716 2904 46722 2916
rect 50338 2904 50344 2916
rect 46716 2876 50344 2904
rect 46716 2864 46722 2876
rect 50338 2864 50344 2876
rect 50396 2864 50402 2916
rect 78582 2864 78588 2916
rect 78640 2904 78646 2916
rect 87248 2904 87276 2944
rect 89162 2932 89168 2984
rect 89220 2972 89226 2984
rect 97258 2972 97264 2984
rect 89220 2944 97264 2972
rect 89220 2932 89226 2944
rect 97258 2932 97264 2944
rect 97316 2932 97322 2984
rect 99834 2932 99840 2984
rect 99892 2972 99898 2984
rect 206278 2972 206284 2984
rect 99892 2944 206284 2972
rect 99892 2932 99898 2944
rect 206278 2932 206284 2944
rect 206336 2932 206342 2984
rect 267734 2932 267740 2984
rect 267792 2972 267798 2984
rect 271138 2972 271144 2984
rect 267792 2944 271144 2972
rect 267792 2932 267798 2944
rect 271138 2932 271144 2944
rect 271196 2932 271202 2984
rect 297266 2932 297272 2984
rect 297324 2972 297330 2984
rect 298370 2972 298376 2984
rect 297324 2944 298376 2972
rect 297324 2932 297330 2944
rect 298370 2932 298376 2944
rect 298428 2932 298434 2984
rect 300762 2932 300768 2984
rect 300820 2972 300826 2984
rect 302237 2975 302295 2981
rect 302237 2972 302249 2975
rect 300820 2944 302249 2972
rect 300820 2932 300826 2944
rect 302237 2941 302249 2944
rect 302283 2941 302295 2975
rect 302344 2972 302372 3012
rect 314010 3000 314016 3012
rect 314068 3000 314074 3052
rect 315022 3000 315028 3052
rect 315080 3040 315086 3052
rect 318058 3040 318064 3052
rect 315080 3012 318064 3040
rect 315080 3000 315086 3012
rect 318058 3000 318064 3012
rect 318116 3000 318122 3052
rect 325666 3040 325694 3080
rect 326709 3077 326721 3111
rect 326755 3108 326767 3111
rect 334158 3108 334164 3120
rect 326755 3080 334164 3108
rect 326755 3077 326767 3080
rect 326709 3071 326767 3077
rect 334158 3068 334164 3080
rect 334216 3068 334222 3120
rect 361114 3068 361120 3120
rect 361172 3108 361178 3120
rect 361172 3080 415440 3108
rect 361172 3068 361178 3080
rect 335998 3040 336004 3052
rect 325666 3012 336004 3040
rect 335998 3000 336004 3012
rect 336056 3000 336062 3052
rect 336274 3000 336280 3052
rect 336332 3040 336338 3052
rect 360838 3040 360844 3052
rect 336332 3012 360844 3040
rect 336332 3000 336338 3012
rect 360838 3000 360844 3012
rect 360896 3000 360902 3052
rect 362310 3000 362316 3052
rect 362368 3040 362374 3052
rect 364978 3040 364984 3052
rect 362368 3012 364984 3040
rect 362368 3000 362374 3012
rect 364978 3000 364984 3012
rect 365036 3000 365042 3052
rect 365806 3000 365812 3052
rect 365864 3040 365870 3052
rect 415305 3043 415363 3049
rect 415305 3040 415317 3043
rect 365864 3012 415317 3040
rect 365864 3000 365870 3012
rect 415305 3009 415317 3012
rect 415351 3009 415363 3043
rect 415412 3040 415440 3080
rect 415486 3068 415492 3120
rect 415544 3108 415550 3120
rect 419537 3111 419595 3117
rect 419537 3108 419549 3111
rect 415544 3080 419549 3108
rect 415544 3068 415550 3080
rect 419537 3077 419549 3080
rect 419583 3077 419595 3111
rect 419537 3071 419595 3077
rect 422570 3068 422576 3120
rect 422628 3108 422634 3120
rect 464338 3108 464344 3120
rect 422628 3080 464344 3108
rect 422628 3068 422634 3080
rect 464338 3068 464344 3080
rect 464396 3068 464402 3120
rect 573910 3068 573916 3120
rect 573968 3108 573974 3120
rect 575566 3108 575572 3120
rect 573968 3080 575572 3108
rect 573968 3068 573974 3080
rect 575566 3068 575572 3080
rect 575624 3068 575630 3120
rect 420086 3040 420092 3052
rect 415412 3012 420092 3040
rect 415305 3003 415363 3009
rect 420086 3000 420092 3012
rect 420144 3000 420150 3052
rect 428458 3000 428464 3052
rect 428516 3040 428522 3052
rect 428516 3012 442580 3040
rect 428516 3000 428522 3012
rect 316678 2972 316684 2984
rect 302344 2944 316684 2972
rect 302237 2935 302295 2941
rect 316678 2932 316684 2944
rect 316736 2932 316742 2984
rect 332686 2932 332692 2984
rect 332744 2972 332750 2984
rect 346854 2972 346860 2984
rect 332744 2944 346860 2972
rect 332744 2932 332750 2944
rect 346854 2932 346860 2944
rect 346912 2932 346918 2984
rect 346946 2932 346952 2984
rect 347004 2972 347010 2984
rect 355321 2975 355379 2981
rect 355321 2972 355333 2975
rect 347004 2944 355333 2972
rect 347004 2932 347010 2944
rect 355321 2941 355333 2944
rect 355367 2941 355379 2975
rect 355321 2935 355379 2941
rect 372890 2932 372896 2984
rect 372948 2972 372954 2984
rect 425698 2972 425704 2984
rect 372948 2944 425704 2972
rect 372948 2932 372954 2944
rect 425698 2932 425704 2944
rect 425756 2932 425762 2984
rect 426158 2932 426164 2984
rect 426216 2972 426222 2984
rect 433153 2975 433211 2981
rect 433153 2972 433165 2975
rect 426216 2944 433165 2972
rect 426216 2932 426222 2944
rect 433153 2941 433165 2944
rect 433199 2941 433211 2975
rect 433153 2935 433211 2941
rect 433242 2932 433248 2984
rect 433300 2972 433306 2984
rect 435453 2975 435511 2981
rect 435453 2972 435465 2975
rect 433300 2944 435465 2972
rect 433300 2932 433306 2944
rect 435453 2941 435465 2944
rect 435499 2941 435511 2975
rect 435453 2935 435511 2941
rect 435542 2932 435548 2984
rect 435600 2972 435606 2984
rect 440237 2975 440295 2981
rect 440237 2972 440249 2975
rect 435600 2944 440249 2972
rect 435600 2932 435606 2944
rect 440237 2941 440249 2944
rect 440283 2941 440295 2975
rect 440237 2935 440295 2941
rect 90266 2904 90272 2916
rect 78640 2876 84194 2904
rect 87248 2876 90272 2904
rect 78640 2864 78646 2876
rect 84166 2836 84194 2876
rect 90266 2864 90272 2876
rect 90324 2864 90330 2916
rect 92750 2864 92756 2916
rect 92808 2904 92814 2916
rect 93302 2904 93308 2916
rect 92808 2876 93308 2904
rect 92808 2864 92814 2876
rect 93302 2864 93308 2876
rect 93360 2864 93366 2916
rect 96246 2864 96252 2916
rect 96304 2904 96310 2916
rect 101398 2904 101404 2916
rect 96304 2876 101404 2904
rect 96304 2864 96310 2876
rect 101398 2864 101404 2876
rect 101456 2864 101462 2916
rect 103330 2864 103336 2916
rect 103388 2904 103394 2916
rect 103388 2876 103514 2904
rect 103388 2864 103394 2876
rect 94498 2836 94504 2848
rect 84166 2808 94504 2836
rect 94498 2796 94504 2808
rect 94556 2796 94562 2848
rect 103486 2836 103514 2876
rect 106918 2864 106924 2916
rect 106976 2904 106982 2916
rect 118697 2907 118755 2913
rect 118697 2904 118709 2907
rect 106976 2876 118709 2904
rect 106976 2864 106982 2876
rect 118697 2873 118709 2876
rect 118743 2873 118755 2907
rect 221642 2904 221648 2916
rect 118697 2867 118755 2873
rect 122806 2876 221648 2904
rect 108298 2836 108304 2848
rect 103486 2808 108304 2836
rect 108298 2796 108304 2808
rect 108356 2796 108362 2848
rect 121086 2796 121092 2848
rect 121144 2836 121150 2848
rect 122806 2836 122834 2876
rect 221642 2864 221648 2876
rect 221700 2864 221706 2916
rect 301958 2864 301964 2916
rect 302016 2904 302022 2916
rect 379698 2904 379704 2916
rect 302016 2876 379704 2904
rect 302016 2864 302022 2876
rect 379698 2864 379704 2876
rect 379756 2864 379762 2916
rect 379974 2864 379980 2916
rect 380032 2904 380038 2916
rect 383013 2907 383071 2913
rect 383013 2904 383025 2907
rect 380032 2876 383025 2904
rect 380032 2864 380038 2876
rect 383013 2873 383025 2876
rect 383059 2873 383071 2907
rect 383013 2867 383071 2873
rect 387150 2864 387156 2916
rect 387208 2904 387214 2916
rect 392673 2907 392731 2913
rect 392673 2904 392685 2907
rect 387208 2876 392685 2904
rect 387208 2864 387214 2876
rect 392673 2873 392685 2876
rect 392719 2873 392731 2907
rect 392673 2867 392731 2873
rect 394234 2864 394240 2916
rect 394292 2904 394298 2916
rect 442258 2904 442264 2916
rect 394292 2876 442264 2904
rect 394292 2864 394298 2876
rect 442258 2864 442264 2876
rect 442316 2864 442322 2916
rect 442552 2904 442580 3012
rect 442626 3000 442632 3052
rect 442684 3040 442690 3052
rect 447778 3040 447784 3052
rect 442684 3012 447784 3040
rect 442684 3000 442690 3012
rect 447778 3000 447784 3012
rect 447836 3000 447842 3052
rect 454494 3000 454500 3052
rect 454552 3040 454558 3052
rect 465721 3043 465779 3049
rect 465721 3040 465733 3043
rect 454552 3012 465733 3040
rect 454552 3000 454558 3012
rect 465721 3009 465733 3012
rect 465767 3009 465779 3043
rect 465721 3003 465779 3009
rect 475746 3000 475752 3052
rect 475804 3040 475810 3052
rect 479610 3040 479616 3052
rect 475804 3012 479616 3040
rect 475804 3000 475810 3012
rect 479610 3000 479616 3012
rect 479668 3000 479674 3052
rect 547874 3000 547880 3052
rect 547932 3040 547938 3052
rect 555418 3040 555424 3052
rect 547932 3012 555424 3040
rect 547932 3000 547938 3012
rect 555418 3000 555424 3012
rect 555476 3000 555482 3052
rect 558546 3000 558552 3052
rect 558604 3040 558610 3052
rect 564618 3040 564624 3052
rect 558604 3012 564624 3040
rect 558604 3000 558610 3012
rect 564618 3000 564624 3012
rect 564676 3000 564682 3052
rect 578602 3000 578608 3052
rect 578660 3040 578666 3052
rect 579614 3040 579620 3052
rect 578660 3012 579620 3040
rect 578660 3000 578666 3012
rect 579614 3000 579620 3012
rect 579672 3000 579678 3052
rect 445018 2932 445024 2984
rect 445076 2972 445082 2984
rect 445754 2972 445760 2984
rect 445076 2944 445760 2972
rect 445076 2932 445082 2944
rect 445754 2932 445760 2944
rect 445812 2932 445818 2984
rect 489914 2932 489920 2984
rect 489972 2972 489978 2984
rect 497458 2972 497464 2984
rect 489972 2944 497464 2972
rect 489972 2932 489978 2944
rect 497458 2932 497464 2944
rect 497516 2932 497522 2984
rect 525426 2932 525432 2984
rect 525484 2972 525490 2984
rect 526438 2972 526444 2984
rect 525484 2944 526444 2972
rect 525484 2932 525490 2944
rect 526438 2932 526444 2944
rect 526496 2932 526502 2984
rect 572714 2932 572720 2984
rect 572772 2972 572778 2984
rect 574186 2972 574192 2984
rect 572772 2944 574192 2972
rect 572772 2932 572778 2944
rect 574186 2932 574192 2944
rect 574244 2932 574250 2984
rect 449158 2904 449164 2916
rect 442552 2876 449164 2904
rect 449158 2864 449164 2876
rect 449216 2864 449222 2916
rect 121144 2808 122834 2836
rect 121144 2796 121150 2808
rect 123478 2796 123484 2848
rect 123536 2836 123542 2848
rect 124122 2836 124128 2848
rect 123536 2808 124128 2836
rect 123536 2796 123542 2808
rect 124122 2796 124128 2808
rect 124180 2796 124186 2848
rect 124674 2796 124680 2848
rect 124732 2836 124738 2848
rect 125410 2836 125416 2848
rect 124732 2808 125416 2836
rect 124732 2796 124738 2808
rect 125410 2796 125416 2808
rect 125468 2796 125474 2848
rect 125870 2796 125876 2848
rect 125928 2836 125934 2848
rect 126882 2836 126888 2848
rect 125928 2808 126888 2836
rect 125928 2796 125934 2808
rect 126882 2796 126888 2808
rect 126940 2796 126946 2848
rect 132954 2796 132960 2848
rect 133012 2836 133018 2848
rect 133782 2836 133788 2848
rect 133012 2808 133788 2836
rect 133012 2796 133018 2808
rect 133782 2796 133788 2808
rect 133840 2796 133846 2848
rect 134150 2796 134156 2848
rect 134208 2836 134214 2848
rect 135162 2836 135168 2848
rect 134208 2808 135168 2836
rect 134208 2796 134214 2808
rect 135162 2796 135168 2808
rect 135220 2796 135226 2848
rect 140038 2796 140044 2848
rect 140096 2836 140102 2848
rect 140682 2836 140688 2848
rect 140096 2808 140688 2836
rect 140096 2796 140102 2808
rect 140682 2796 140688 2808
rect 140740 2796 140746 2848
rect 141234 2796 141240 2848
rect 141292 2836 141298 2848
rect 142062 2836 142068 2848
rect 141292 2808 142068 2836
rect 141292 2796 141298 2808
rect 142062 2796 142068 2808
rect 142120 2796 142126 2848
rect 143534 2796 143540 2848
rect 143592 2836 143598 2848
rect 144822 2836 144828 2848
rect 143592 2808 144828 2836
rect 143592 2796 143598 2808
rect 144822 2796 144828 2808
rect 144880 2796 144886 2848
rect 147122 2796 147128 2848
rect 147180 2836 147186 2848
rect 147582 2836 147588 2848
rect 147180 2808 147588 2836
rect 147180 2796 147186 2808
rect 147582 2796 147588 2808
rect 147640 2796 147646 2848
rect 148318 2796 148324 2848
rect 148376 2836 148382 2848
rect 148962 2836 148968 2848
rect 148376 2808 148968 2836
rect 148376 2796 148382 2808
rect 148962 2796 148968 2808
rect 149020 2796 149026 2848
rect 150618 2796 150624 2848
rect 150676 2836 150682 2848
rect 151722 2836 151728 2848
rect 150676 2808 151728 2836
rect 150676 2796 150682 2808
rect 151722 2796 151728 2808
rect 151780 2796 151786 2848
rect 151814 2796 151820 2848
rect 151872 2836 151878 2848
rect 153102 2836 153108 2848
rect 151872 2808 153108 2836
rect 151872 2796 151878 2808
rect 153102 2796 153108 2808
rect 153160 2796 153166 2848
rect 155402 2796 155408 2848
rect 155460 2836 155466 2848
rect 155862 2836 155868 2848
rect 155460 2808 155868 2836
rect 155460 2796 155466 2808
rect 155862 2796 155868 2808
rect 155920 2796 155926 2848
rect 157794 2796 157800 2848
rect 157852 2836 157858 2848
rect 158622 2836 158628 2848
rect 157852 2808 158628 2836
rect 157852 2796 157858 2808
rect 158622 2796 158628 2808
rect 158680 2796 158686 2848
rect 158898 2796 158904 2848
rect 158956 2836 158962 2848
rect 160002 2836 160008 2848
rect 158956 2808 160008 2836
rect 158956 2796 158962 2808
rect 160002 2796 160008 2808
rect 160060 2796 160066 2848
rect 164789 2839 164847 2845
rect 164789 2805 164801 2839
rect 164835 2836 164847 2839
rect 169846 2836 169852 2848
rect 164835 2808 169852 2836
rect 164835 2805 164847 2808
rect 164789 2799 164847 2805
rect 169846 2796 169852 2808
rect 169904 2796 169910 2848
rect 298281 2839 298339 2845
rect 298281 2805 298293 2839
rect 298327 2836 298339 2839
rect 302878 2836 302884 2848
rect 298327 2808 302884 2836
rect 298327 2805 298339 2808
rect 298281 2799 298339 2805
rect 302878 2796 302884 2808
rect 302936 2796 302942 2848
rect 396534 2796 396540 2848
rect 396592 2836 396598 2848
rect 399573 2839 399631 2845
rect 399573 2836 399585 2839
rect 396592 2808 399585 2836
rect 396592 2796 396598 2808
rect 399573 2805 399585 2808
rect 399619 2805 399631 2839
rect 399573 2799 399631 2805
rect 404725 2839 404783 2845
rect 404725 2805 404737 2839
rect 404771 2836 404783 2839
rect 412726 2836 412732 2848
rect 404771 2808 412732 2836
rect 404771 2805 404783 2808
rect 404725 2799 404783 2805
rect 412726 2796 412732 2808
rect 412784 2796 412790 2848
rect 417878 2796 417884 2848
rect 417936 2836 417942 2848
rect 454678 2836 454684 2848
rect 417936 2808 454684 2836
rect 417936 2796 417942 2808
rect 454678 2796 454684 2808
rect 454736 2796 454742 2848
<< via1 >>
rect 141424 703604 141476 703656
rect 551100 703604 551152 703656
rect 345020 703536 345072 703588
rect 396356 703536 396408 703588
rect 342168 703468 342220 703520
rect 407396 703468 407448 703520
rect 275468 703400 275520 703452
rect 351184 703400 351236 703452
rect 352840 703400 352892 703452
rect 429844 703400 429896 703452
rect 161572 703332 161624 703384
rect 346400 703332 346452 703384
rect 349068 703332 349120 703384
rect 478512 703332 478564 703384
rect 235172 703264 235224 703316
rect 385316 703264 385368 703316
rect 340420 703196 340472 703248
rect 577044 703196 577096 703248
rect 164792 703128 164844 703180
rect 440608 703128 440660 703180
rect 164516 703060 164568 703112
rect 451648 703060 451700 703112
rect 282828 702992 282880 703044
rect 576952 702992 577004 703044
rect 165344 702924 165396 702976
rect 462688 702924 462740 702976
rect 165160 702856 165212 702908
rect 473728 702856 473780 702908
rect 161848 702788 161900 702840
rect 484768 702788 484820 702840
rect 162032 702720 162084 702772
rect 495808 702720 495860 702772
rect 231216 702652 231268 702704
rect 198096 702584 198148 702636
rect 148324 702516 148376 702568
rect 540060 702516 540112 702568
rect 356060 702448 356112 702500
rect 374276 702448 374328 702500
rect 14464 702380 14516 702432
rect 466460 702380 466512 702432
rect 17224 702312 17276 702364
rect 477500 702312 477552 702364
rect 341800 702244 341852 702296
rect 350448 702244 350500 702296
rect 351184 702244 351236 702296
rect 362500 702244 362552 702296
rect 363880 702244 363932 702296
rect 364984 702244 365036 702296
rect 367192 702287 367244 702296
rect 367192 702253 367201 702287
rect 367201 702253 367235 702287
rect 367235 702253 367244 702287
rect 367192 702244 367244 702253
rect 323308 702176 323360 702228
rect 419356 702176 419408 702228
rect 253388 702108 253440 702160
rect 340420 702108 340472 702160
rect 346400 702108 346452 702160
rect 447968 702108 448020 702160
rect 71044 702040 71096 702092
rect 358728 702040 358780 702092
rect 65524 701972 65576 702024
rect 360292 702040 360344 702092
rect 359096 701972 359148 702024
rect 392676 702040 392728 702092
rect 361764 701972 361816 702024
rect 547420 701972 547472 702024
rect 293546 701904 293598 701956
rect 583484 701904 583536 701956
rect 289866 701836 289918 701888
rect 583576 701836 583628 701888
rect 161664 701768 161716 701820
rect 459008 701768 459060 701820
rect 562784 701768 562836 701820
rect 279148 701700 279200 701752
rect 583392 701700 583444 701752
rect 161756 701632 161808 701684
rect 470048 701632 470100 701684
rect 555424 701632 555476 701684
rect 162124 701564 162176 701616
rect 161940 701496 161992 701548
rect 271788 701564 271840 701616
rect 583208 701564 583260 701616
rect 162400 701428 162452 701480
rect 162216 701360 162268 701412
rect 179052 701496 179104 701548
rect 268108 701496 268160 701548
rect 583300 701496 583352 701548
rect 190092 701428 190144 701480
rect 260748 701428 260800 701480
rect 583024 701428 583076 701480
rect 162492 701292 162544 701344
rect 162308 701224 162360 701276
rect 492128 701360 492180 701412
rect 566464 701360 566516 701412
rect 182732 701292 182784 701344
rect 249708 701292 249760 701344
rect 582840 701292 582892 701344
rect 162584 701156 162636 701208
rect 168012 701156 168064 701208
rect 186412 701224 186464 701276
rect 245752 701224 245804 701276
rect 582932 701224 582984 701276
rect 162768 701088 162820 701140
rect 164332 701088 164384 701140
rect 170312 701131 170364 701140
rect 170312 701097 170321 701131
rect 170321 701097 170355 701131
rect 170355 701097 170364 701131
rect 170312 701088 170364 701097
rect 162676 701020 162728 701072
rect 171692 701156 171744 701208
rect 242256 701156 242308 701208
rect 583760 701156 583812 701208
rect 175372 701088 175424 701140
rect 202788 701131 202840 701140
rect 202788 701097 202797 701131
rect 202797 701097 202831 701131
rect 202831 701097 202840 701131
rect 202788 701088 202840 701097
rect 257068 701131 257120 701140
rect 257068 701097 257077 701131
rect 257077 701097 257111 701131
rect 257111 701097 257120 701131
rect 257068 701088 257120 701097
rect 267648 701131 267700 701140
rect 267648 701097 267657 701131
rect 267657 701097 267691 701131
rect 267691 701097 267700 701131
rect 267648 701088 267700 701097
rect 283840 701131 283892 701140
rect 283840 701097 283849 701131
rect 283849 701097 283883 701131
rect 283883 701097 283892 701131
rect 283840 701088 283892 701097
rect 300124 701131 300176 701140
rect 300124 701097 300133 701131
rect 300133 701097 300167 701131
rect 300167 701097 300176 701131
rect 300124 701088 300176 701097
rect 304908 701131 304960 701140
rect 304908 701097 304917 701131
rect 304917 701097 304951 701131
rect 304951 701097 304960 701131
rect 304908 701088 304960 701097
rect 330208 701131 330260 701140
rect 330208 701097 330217 701131
rect 330217 701097 330251 701131
rect 330251 701097 330260 701131
rect 330208 701088 330260 701097
rect 332508 701131 332560 701140
rect 332508 701097 332517 701131
rect 332517 701097 332551 701131
rect 332551 701097 332560 701131
rect 332508 701088 332560 701097
rect 338028 701088 338080 701140
rect 342168 701131 342220 701140
rect 342168 701097 342177 701131
rect 342177 701097 342211 701131
rect 342211 701097 342220 701131
rect 342168 701088 342220 701097
rect 345020 701131 345072 701140
rect 345020 701097 345029 701131
rect 345029 701097 345063 701131
rect 345063 701097 345072 701131
rect 345480 701131 345532 701140
rect 345020 701088 345072 701097
rect 345480 701097 345489 701131
rect 345489 701097 345523 701131
rect 345523 701097 345532 701131
rect 345480 701088 345532 701097
rect 348700 701131 348752 701140
rect 348700 701097 348709 701131
rect 348709 701097 348743 701131
rect 348743 701097 348752 701131
rect 348700 701088 348752 701097
rect 356060 701088 356112 701140
rect 356520 701131 356572 701140
rect 356520 701097 356529 701131
rect 356529 701097 356563 701131
rect 356563 701097 356572 701131
rect 356520 701088 356572 701097
rect 359464 701088 359516 701140
rect 367100 701088 367152 701140
rect 370596 701088 370648 701140
rect 378140 701131 378192 701140
rect 378140 701097 378149 701131
rect 378149 701097 378183 701131
rect 378183 701097 378192 701131
rect 378140 701088 378192 701097
rect 381636 701131 381688 701140
rect 381636 701097 381645 701131
rect 381645 701097 381679 701131
rect 381679 701097 381688 701131
rect 381636 701088 381688 701097
rect 389180 701131 389232 701140
rect 389180 701097 389189 701131
rect 389189 701097 389223 701131
rect 389223 701097 389232 701131
rect 389180 701088 389232 701097
rect 397460 701131 397512 701140
rect 397460 701097 397469 701131
rect 397469 701097 397503 701131
rect 397503 701097 397512 701131
rect 397460 701088 397512 701097
rect 400220 701088 400272 701140
rect 403716 701131 403768 701140
rect 403716 701097 403725 701131
rect 403725 701097 403759 701131
rect 403759 701097 403768 701131
rect 403716 701088 403768 701097
rect 411260 701131 411312 701140
rect 411260 701097 411269 701131
rect 411269 701097 411303 701131
rect 411303 701097 411312 701131
rect 411260 701088 411312 701097
rect 413652 701088 413704 701140
rect 414756 701131 414808 701140
rect 414756 701097 414765 701131
rect 414765 701097 414799 701131
rect 414799 701097 414808 701131
rect 414756 701088 414808 701097
rect 422392 701131 422444 701140
rect 422392 701097 422401 701131
rect 422401 701097 422435 701131
rect 422435 701097 422444 701131
rect 422392 701088 422444 701097
rect 425888 701131 425940 701140
rect 425888 701097 425897 701131
rect 425897 701097 425931 701131
rect 425931 701097 425940 701131
rect 425888 701088 425940 701097
rect 433340 701131 433392 701140
rect 433340 701097 433349 701131
rect 433349 701097 433383 701131
rect 433383 701097 433392 701131
rect 433340 701088 433392 701097
rect 436928 701131 436980 701140
rect 436928 701097 436937 701131
rect 436937 701097 436971 701131
rect 436971 701097 436980 701131
rect 436928 701088 436980 701097
rect 444380 701131 444432 701140
rect 444380 701097 444389 701131
rect 444389 701097 444423 701131
rect 444423 701097 444432 701131
rect 444380 701088 444432 701097
rect 455420 701131 455472 701140
rect 455420 701097 455429 701131
rect 455429 701097 455463 701131
rect 455463 701097 455472 701131
rect 455420 701088 455472 701097
rect 462320 701131 462372 701140
rect 462320 701097 462329 701131
rect 462329 701097 462363 701131
rect 462363 701097 462372 701131
rect 462320 701088 462372 701097
rect 543464 701088 543516 701140
rect 543740 701088 543792 701140
rect 558460 701088 558512 701140
rect 569960 701088 570012 701140
rect 137836 700952 137888 701004
rect 105452 700884 105504 700936
rect 53104 700476 53156 700528
rect 154120 700408 154172 700460
rect 3424 700340 3476 700392
rect 577504 701088 577556 701140
rect 583668 700272 583720 700324
rect 583116 700204 583168 700256
rect 89168 700136 89220 700188
rect 72976 700068 73028 700120
rect 35164 700000 35216 700052
rect 24308 699932 24360 699984
rect 40684 699864 40736 699916
rect 43444 699796 43496 699848
rect 8116 699728 8168 699780
rect 14556 699660 14608 699712
rect 3056 671984 3108 672036
rect 35164 671984 35216 672036
rect 3516 658180 3568 658232
rect 14556 658180 14608 658232
rect 3332 619556 3384 619608
rect 161572 619556 161624 619608
rect 3240 607112 3292 607164
rect 40684 607112 40736 607164
rect 3516 567128 3568 567180
rect 161664 567128 161716 567180
rect 3516 554684 3568 554736
rect 43444 554684 43496 554736
rect 3516 516060 3568 516112
rect 161756 516060 161808 516112
rect 3516 502256 3568 502308
rect 14464 502256 14516 502308
rect 3240 463632 3292 463684
rect 32404 463632 32456 463684
rect 3332 449828 3384 449880
rect 17224 449828 17276 449880
rect 3516 423580 3568 423632
rect 161848 423580 161900 423632
rect 2964 411204 3016 411256
rect 161940 411204 161992 411256
rect 3240 398760 3292 398812
rect 18604 398760 18656 398812
rect 3516 372512 3568 372564
rect 162032 372512 162084 372564
rect 3148 346332 3200 346384
rect 79324 346332 79376 346384
rect 3424 306280 3476 306332
rect 29644 306280 29696 306332
rect 3056 293904 3108 293956
rect 105544 293904 105596 293956
rect 162308 282276 162360 282328
rect 580264 282276 580316 282328
rect 162124 282208 162176 282260
rect 580356 282208 580408 282260
rect 162216 282140 162268 282192
rect 580448 282140 580500 282192
rect 97264 280100 97316 280152
rect 226708 280100 226760 280152
rect 226984 280100 227036 280152
rect 246304 280100 246356 280152
rect 320088 280100 320140 280152
rect 351920 280100 351972 280152
rect 352564 280100 352616 280152
rect 414940 280100 414992 280152
rect 419448 280100 419500 280152
rect 464344 280100 464396 280152
rect 471888 280100 471940 280152
rect 501880 280100 501932 280152
rect 503628 280100 503680 280152
rect 524880 280100 524932 280152
rect 525156 280100 525208 280152
rect 540244 280100 540296 280152
rect 576860 280100 576912 280152
rect 577688 280100 577740 280152
rect 111708 280032 111760 280084
rect 242072 280032 242124 280084
rect 255412 280032 255464 280084
rect 261668 280032 261720 280084
rect 302884 280032 302936 280084
rect 367284 280032 367336 280084
rect 369768 280032 369820 280084
rect 428648 280032 428700 280084
rect 430488 280032 430540 280084
rect 472072 280032 472124 280084
rect 472624 280032 472676 280084
rect 484860 280032 484912 280084
rect 485688 280032 485740 280084
rect 512092 280032 512144 280084
rect 513288 280032 513340 280084
rect 531688 280032 531740 280084
rect 533436 280032 533488 280084
rect 545304 280032 545356 280084
rect 101404 279964 101456 280016
rect 231860 279964 231912 280016
rect 295984 279964 296036 280016
rect 313556 279964 313608 280016
rect 323860 279964 323912 280016
rect 35164 279896 35216 279948
rect 179880 279896 179932 279948
rect 222844 279896 222896 279948
rect 248880 279896 248932 279948
rect 249064 279896 249116 279948
rect 260840 279896 260892 279948
rect 276664 279896 276716 279948
rect 318800 279896 318852 279948
rect 322204 279896 322256 279948
rect 325792 279964 325844 280016
rect 326344 279964 326396 280016
rect 328920 279964 328972 280016
rect 329104 279964 329156 280016
rect 397920 279964 397972 280016
rect 399484 279964 399536 280016
rect 449072 279964 449124 280016
rect 449808 279964 449860 280016
rect 486516 279964 486568 280016
rect 496728 279964 496780 280016
rect 519728 279964 519780 280016
rect 527456 279964 527508 280016
rect 537668 279964 537720 280016
rect 538128 279964 538180 280016
rect 549536 279964 549588 280016
rect 392860 279896 392912 279948
rect 393964 279896 394016 279948
rect 50344 279828 50396 279880
rect 196072 279828 196124 279880
rect 196624 279828 196676 279880
rect 216680 279828 216732 279880
rect 221464 279828 221516 279880
rect 43444 279760 43496 279812
rect 190920 279760 190972 279812
rect 199384 279760 199436 279812
rect 221556 279760 221608 279812
rect 221740 279828 221792 279880
rect 249800 279828 249852 279880
rect 252008 279828 252060 279880
rect 278780 279828 278832 279880
rect 309140 279828 309192 279880
rect 310152 279828 310204 279880
rect 313188 279828 313240 279880
rect 387800 279828 387852 279880
rect 244556 279760 244608 279812
rect 244924 279760 244976 279812
rect 283748 279760 283800 279812
rect 306288 279760 306340 279812
rect 382556 279760 382608 279812
rect 384396 279760 384448 279812
rect 389824 279760 389876 279812
rect 390560 279760 390612 279812
rect 394700 279828 394752 279880
rect 395344 279828 395396 279880
rect 400128 279896 400180 279948
rect 450728 279896 450780 279948
rect 454684 279896 454736 279948
rect 463700 279896 463752 279948
rect 466368 279896 466420 279948
rect 497648 279896 497700 279948
rect 502248 279896 502300 279948
rect 524052 279896 524104 279948
rect 525064 279896 525116 279948
rect 539600 279896 539652 279948
rect 543004 279896 543056 279948
rect 552940 279896 552992 279948
rect 445760 279828 445812 279880
rect 451188 279828 451240 279880
rect 487344 279828 487396 279880
rect 489828 279828 489880 279880
rect 514760 279828 514812 279880
rect 516048 279828 516100 279880
rect 534264 279828 534316 279880
rect 536748 279828 536800 279880
rect 548708 279828 548760 279880
rect 438860 279760 438912 279812
rect 440148 279760 440200 279812
rect 478880 279760 478932 279812
rect 482928 279760 482980 279812
rect 509516 279760 509568 279812
rect 514668 279760 514720 279812
rect 532700 279760 532752 279812
rect 533344 279760 533396 279812
rect 546132 279760 546184 279812
rect 547144 279760 547196 279812
rect 555516 279760 555568 279812
rect 36544 279692 36596 279744
rect 185860 279692 185912 279744
rect 208492 279692 208544 279744
rect 251456 279692 251508 279744
rect 251824 279692 251876 279744
rect 254860 279692 254912 279744
rect 281540 279692 281592 279744
rect 299388 279692 299440 279744
rect 377496 279692 377548 279744
rect 377588 279692 377640 279744
rect 433708 279692 433760 279744
rect 437388 279692 437440 279744
rect 477132 279692 477184 279744
rect 479524 279692 479576 279744
rect 506940 279692 506992 279744
rect 507768 279692 507820 279744
rect 519544 279692 519596 279744
rect 526536 279692 526588 279744
rect 535368 279692 535420 279744
rect 548064 279692 548116 279744
rect 549168 279692 549220 279744
rect 558092 279692 558144 279744
rect 29644 279624 29696 279676
rect 180892 279624 180944 279676
rect 187700 279624 187752 279676
rect 188344 279624 188396 279676
rect 200764 279624 200816 279676
rect 224132 279624 224184 279676
rect 233884 279624 233936 279676
rect 286324 279624 286376 279676
rect 293224 279624 293276 279676
rect 372620 279624 372672 279676
rect 373264 279624 373316 279676
rect 425704 279624 425756 279676
rect 431132 279624 431184 279676
rect 433248 279624 433300 279676
rect 473728 279624 473780 279676
rect 480904 279624 480956 279676
rect 507860 279624 507912 279676
rect 509148 279624 509200 279676
rect 529112 279624 529164 279676
rect 529848 279624 529900 279676
rect 543740 279624 543792 279676
rect 544384 279624 544436 279676
rect 553860 279624 553912 279676
rect 558184 279624 558236 279676
rect 562324 279624 562376 279676
rect 572720 279624 572772 279676
rect 573456 279624 573508 279676
rect 582288 279624 582340 279676
rect 18604 279556 18656 279608
rect 173072 279556 173124 279608
rect 195244 279556 195296 279608
rect 211344 279556 211396 279608
rect 214564 279556 214616 279608
rect 239496 279556 239548 279608
rect 242808 279556 242860 279608
rect 317512 279556 317564 279608
rect 321560 279556 321612 279608
rect 327080 279556 327132 279608
rect 328092 279556 328144 279608
rect 334072 279556 334124 279608
rect 334900 279556 334952 279608
rect 403164 279556 403216 279608
rect 407764 279556 407816 279608
rect 410708 279556 410760 279608
rect 454132 279556 454184 279608
rect 458088 279556 458140 279608
rect 492680 279556 492732 279608
rect 493324 279556 493376 279608
rect 517520 279556 517572 279608
rect 522948 279556 523000 279608
rect 538496 279556 538548 279608
rect 539508 279556 539560 279608
rect 550640 279556 550692 279608
rect 558276 279556 558328 279608
rect 563244 279556 563296 279608
rect 572628 279556 572680 279608
rect 574284 279556 574336 279608
rect 17224 279488 17276 279540
rect 173900 279488 173952 279540
rect 191104 279488 191156 279540
rect 201132 279488 201184 279540
rect 203524 279488 203576 279540
rect 229376 279488 229428 279540
rect 251916 279488 251968 279540
rect 341708 279488 341760 279540
rect 342904 279488 342956 279540
rect 344284 279488 344336 279540
rect 349068 279488 349120 279540
rect 413284 279488 413336 279540
rect 415308 279488 415360 279540
rect 461032 279488 461084 279540
rect 464436 279488 464488 279540
rect 466092 279488 466144 279540
rect 467104 279488 467156 279540
rect 469496 279488 469548 279540
rect 494152 279488 494204 279540
rect 495348 279488 495400 279540
rect 518900 279488 518952 279540
rect 520188 279488 520240 279540
rect 536840 279488 536892 279540
rect 540888 279488 540940 279540
rect 552112 279488 552164 279540
rect 554688 279488 554740 279540
rect 561680 279488 561732 279540
rect 569224 279488 569276 279540
rect 571708 279488 571760 279540
rect 7564 279420 7616 279472
rect 167092 279420 167144 279472
rect 169760 279420 169812 279472
rect 170496 279420 170548 279472
rect 180064 279420 180116 279472
rect 190092 279420 190144 279472
rect 192484 279420 192536 279472
rect 206284 279420 206336 279472
rect 206376 279420 206428 279472
rect 234620 279420 234672 279472
rect 242716 279420 242768 279472
rect 336740 279420 336792 279472
rect 342168 279420 342220 279472
rect 408132 279420 408184 279472
rect 412548 279420 412600 279472
rect 459560 279420 459612 279472
rect 464344 279420 464396 279472
rect 466920 279420 466972 279472
rect 467748 279420 467800 279472
rect 499580 279420 499632 279472
rect 500868 279420 500920 279472
rect 523132 279420 523184 279472
rect 526444 279420 526496 279472
rect 541072 279420 541124 279472
rect 545028 279420 545080 279472
rect 554780 279420 554832 279472
rect 557448 279420 557500 279472
rect 564072 279420 564124 279472
rect 565728 279420 565780 279472
rect 570052 279420 570104 279472
rect 118608 279352 118660 279404
rect 247132 279352 247184 279404
rect 249708 279352 249760 279404
rect 269120 279352 269172 279404
rect 270132 279352 270184 279404
rect 300124 279352 300176 279404
rect 357072 279352 357124 279404
rect 358820 279352 358872 279404
rect 359556 279352 359608 279404
rect 418344 279352 418396 279404
rect 421564 279352 421616 279404
rect 426072 279352 426124 279404
rect 431224 279352 431276 279404
rect 436284 279352 436336 279404
rect 444288 279352 444340 279404
rect 482284 279352 482336 279404
rect 487068 279352 487120 279404
rect 512920 279352 512972 279404
rect 515956 279352 516008 279404
rect 533528 279352 533580 279404
rect 108304 279284 108356 279336
rect 236920 279284 236972 279336
rect 316040 279284 316092 279336
rect 316960 279284 317012 279336
rect 323584 279284 323636 279336
rect 346860 279284 346912 279336
rect 358728 279284 358780 279336
rect 420092 279284 420144 279336
rect 430580 279284 430632 279336
rect 461584 279284 461636 279336
rect 491668 279284 491720 279336
rect 501604 279284 501656 279336
rect 520648 279284 520700 279336
rect 527088 279284 527140 279336
rect 541900 279284 541952 279336
rect 125508 279216 125560 279268
rect 252560 279216 252612 279268
rect 307024 279216 307076 279268
rect 362132 279216 362184 279268
rect 364984 279216 365036 279268
rect 423680 279216 423732 279268
rect 454776 279216 454828 279268
rect 458456 279216 458508 279268
rect 460296 279216 460348 279268
rect 489092 279216 489144 279268
rect 502984 279216 503036 279268
rect 506112 279216 506164 279268
rect 511908 279216 511960 279268
rect 530860 279216 530912 279268
rect 531228 279216 531280 279268
rect 544476 279216 544528 279268
rect 548524 279216 548576 279268
rect 556344 279216 556396 279268
rect 561588 279216 561640 279268
rect 566648 279216 566700 279268
rect 94504 279148 94556 279200
rect 219072 279148 219124 279200
rect 313924 279148 313976 279200
rect 331496 279148 331548 279200
rect 333888 279148 333940 279200
rect 356704 279148 356756 279200
rect 366364 279148 366416 279200
rect 425152 279148 425204 279200
rect 449164 279148 449216 279200
rect 471152 279148 471204 279200
rect 479616 279148 479668 279200
rect 505284 279148 505336 279200
rect 517428 279148 517480 279200
rect 535092 279148 535144 279200
rect 90364 279080 90416 279132
rect 208860 279080 208912 279132
rect 320824 279080 320876 279132
rect 379428 279080 379480 279132
rect 435456 279080 435508 279132
rect 456064 279080 456116 279132
rect 476304 279080 476356 279132
rect 478144 279080 478196 279132
rect 502708 279080 502760 279132
rect 504364 279080 504416 279132
rect 518072 279080 518124 279132
rect 518164 279080 518216 279132
rect 529940 279080 529992 279132
rect 87604 279012 87656 279064
rect 203708 279012 203760 279064
rect 388444 279012 388496 279064
rect 440516 279012 440568 279064
rect 86224 278944 86276 278996
rect 198740 278944 198792 278996
rect 391848 278944 391900 278996
rect 443920 279012 443972 279064
rect 460204 279012 460256 279064
rect 483940 279012 483992 279064
rect 497464 279012 497516 279064
rect 515496 279012 515548 279064
rect 521568 279012 521620 279064
rect 442264 278944 442316 278996
rect 446496 278944 446548 278996
rect 468484 278944 468536 278996
rect 474740 278944 474792 278996
rect 476764 278944 476816 278996
rect 500132 278944 500184 278996
rect 508504 278944 508556 278996
rect 521660 278944 521712 278996
rect 106924 278876 106976 278928
rect 213920 278876 213972 278928
rect 409144 278876 409196 278928
rect 455880 278876 455932 278928
rect 462964 278876 463016 278928
rect 475384 278876 475436 278928
rect 495072 278876 495124 278928
rect 512644 278876 512696 278928
rect 525800 278876 525852 278928
rect 551284 278876 551336 278928
rect 558920 278876 558972 278928
rect 262312 278808 262364 278860
rect 265900 278808 265952 278860
rect 405648 278808 405700 278860
rect 474004 278808 474056 278860
rect 490012 278808 490064 278860
rect 556804 278808 556856 278860
rect 559748 278808 559800 278860
rect 562968 278808 563020 278860
rect 567476 278808 567528 278860
rect 349804 278740 349856 278792
rect 354680 278740 354732 278792
rect 363604 278740 363656 278792
rect 364708 278740 364760 278792
rect 383016 278740 383068 278792
rect 384304 278740 384356 278792
rect 420184 278740 420236 278792
rect 422668 278740 422720 278792
rect 436744 278740 436796 278792
rect 441620 278740 441672 278792
rect 469864 278740 469916 278792
rect 479708 278740 479760 278792
rect 555424 278740 555476 278792
rect 557540 278740 557592 278792
rect 566464 278740 566516 278792
rect 569132 278740 569184 278792
rect 575388 278740 575440 278792
rect 576952 278740 577004 278792
rect 115204 278672 115256 278724
rect 243728 278672 243780 278724
rect 278044 278672 278096 278724
rect 351092 278672 351144 278724
rect 364248 278672 364300 278724
rect 424232 278672 424284 278724
rect 424324 278672 424376 278724
rect 465264 278672 465316 278724
rect 39304 278604 39356 278656
rect 172152 278604 172204 278656
rect 291844 278604 291896 278656
rect 366456 278604 366508 278656
rect 367744 278604 367796 278656
rect 426900 278604 426952 278656
rect 447784 278604 447836 278656
rect 481640 278604 481692 278656
rect 99288 278536 99340 278588
rect 233148 278536 233200 278588
rect 289084 278536 289136 278588
rect 368940 278536 368992 278588
rect 375288 278536 375340 278588
rect 432052 278536 432104 278588
rect 435364 278536 435416 278588
rect 475476 278536 475528 278588
rect 32404 278468 32456 278520
rect 167920 278468 167972 278520
rect 209044 278468 209096 278520
rect 293960 278468 294012 278520
rect 314016 278468 314068 278520
rect 379152 278468 379204 278520
rect 382924 278468 382976 278520
rect 437112 278468 437164 278520
rect 440884 278468 440936 278520
rect 478052 278468 478104 278520
rect 486424 278468 486476 278520
rect 495900 278536 495952 278588
rect 95056 278400 95108 278452
rect 230940 278400 230992 278452
rect 271144 278400 271196 278452
rect 355324 278400 355376 278452
rect 360108 278400 360160 278452
rect 421748 278400 421800 278452
rect 425796 278400 425848 278452
rect 467840 278400 467892 278452
rect 485044 278400 485096 278452
rect 493508 278468 493560 278520
rect 493416 278400 493468 278452
rect 503720 278400 503772 278452
rect 88984 278332 89036 278384
rect 225880 278332 225932 278384
rect 258724 278332 258776 278384
rect 343640 278332 343692 278384
rect 357348 278332 357400 278384
rect 419540 278332 419592 278384
rect 428464 278332 428516 278384
rect 470600 278332 470652 278384
rect 482284 278332 482336 278384
rect 508688 278332 508740 278384
rect 25504 278264 25556 278316
rect 164516 278264 164568 278316
rect 224868 278264 224920 278316
rect 242808 278264 242860 278316
rect 260104 278264 260156 278316
rect 348516 278264 348568 278316
rect 353944 278264 353996 278316
rect 416780 278264 416832 278316
rect 417424 278264 417476 278316
rect 462688 278264 462740 278316
rect 484308 278264 484360 278316
rect 511264 278264 511316 278316
rect 81348 278196 81400 278248
rect 220820 278196 220872 278248
rect 242164 278196 242216 278248
rect 332600 278196 332652 278248
rect 342076 278196 342128 278248
rect 409052 278196 409104 278248
rect 410524 278196 410576 278248
rect 457536 278196 457588 278248
rect 471244 278196 471296 278248
rect 501052 278196 501104 278248
rect 22744 278128 22796 278180
rect 163688 278128 163740 278180
rect 240784 278128 240836 278180
rect 333152 278128 333204 278180
rect 339408 278128 339460 278180
rect 406476 278128 406528 278180
rect 407028 278128 407080 278180
rect 455052 278128 455104 278180
rect 466276 278128 466328 278180
rect 498476 278128 498528 278180
rect 48228 278060 48280 278112
rect 196900 278060 196952 278112
rect 233148 278060 233200 278112
rect 329840 278060 329892 278112
rect 331864 278060 331916 278112
rect 399668 278060 399720 278112
rect 400864 278060 400916 278112
rect 449900 278060 449952 278112
rect 450544 278060 450596 278112
rect 485780 278060 485832 278112
rect 489184 278060 489236 278112
rect 513748 278060 513800 278112
rect 14464 277992 14516 278044
rect 162860 277992 162912 278044
rect 227628 277992 227680 278044
rect 325884 277992 325936 278044
rect 332508 277992 332560 278044
rect 401600 277992 401652 278044
rect 403624 277992 403676 278044
rect 452660 277992 452712 278044
rect 453304 277992 453356 278044
rect 488540 277992 488592 278044
rect 491208 277992 491260 278044
rect 516324 277992 516376 278044
rect 135168 277924 135220 277976
rect 259092 277924 259144 277976
rect 316684 277924 316736 277976
rect 374092 277924 374144 277976
rect 392584 277924 392636 277976
rect 444748 277924 444800 277976
rect 446404 277924 446456 277976
rect 480536 277924 480588 277976
rect 151728 277856 151780 277908
rect 270960 277856 271012 277908
rect 336004 277856 336056 277908
rect 386880 277856 386932 277908
rect 389916 277856 389968 277908
rect 442356 277856 442408 277908
rect 144828 277788 144880 277840
rect 262312 277788 262364 277840
rect 396724 277788 396776 277840
rect 447324 277788 447376 277840
rect 246304 277720 246356 277772
rect 311900 277720 311952 277772
rect 413928 277720 413980 277772
rect 460112 277720 460164 277772
rect 231124 277652 231176 277704
rect 296720 277652 296772 277704
rect 250444 277584 250496 277636
rect 314660 277584 314712 277636
rect 238024 277516 238076 277568
rect 301688 277516 301740 277568
rect 262864 277448 262916 277500
rect 319536 277448 319588 277500
rect 253204 277380 253256 277432
rect 299112 277380 299164 277432
rect 137928 277312 137980 277364
rect 255412 277312 255464 277364
rect 153108 277244 153160 277296
rect 271788 277244 271840 277296
rect 273904 277244 273956 277296
rect 340972 277244 341024 277296
rect 155868 277176 155920 277228
rect 274548 277176 274600 277228
rect 112444 277108 112496 277160
rect 240232 277108 240284 277160
rect 267004 277108 267056 277160
rect 338212 277108 338264 277160
rect 347044 277108 347096 277160
rect 401784 277108 401836 277160
rect 105544 277040 105596 277092
rect 236092 277040 236144 277092
rect 280804 277040 280856 277092
rect 356152 277040 356204 277092
rect 54484 276972 54536 277024
rect 185032 276972 185084 277024
rect 284944 276972 284996 277024
rect 361580 276972 361632 277024
rect 106188 276904 106240 276956
rect 238668 276904 238720 276956
rect 286324 276904 286376 276956
rect 363052 276904 363104 276956
rect 58624 276836 58676 276888
rect 191932 276836 191984 276888
rect 220728 276836 220780 276888
rect 317512 276836 317564 276888
rect 324964 276836 325016 276888
rect 394792 276836 394844 276888
rect 93124 276768 93176 276820
rect 227996 276768 228048 276820
rect 282184 276768 282236 276820
rect 358912 276768 358964 276820
rect 360844 276768 360896 276820
rect 404360 276768 404412 276820
rect 40684 276700 40736 276752
rect 178132 276700 178184 276752
rect 227536 276700 227588 276752
rect 325608 276700 325660 276752
rect 340144 276700 340196 276752
rect 396172 276700 396224 276752
rect 33784 276632 33836 276684
rect 175280 276632 175332 276684
rect 215944 276632 215996 276684
rect 316132 276632 316184 276684
rect 318064 276632 318116 276684
rect 389180 276632 389232 276684
rect 431868 276632 431920 276684
rect 472072 276632 472124 276684
rect 160008 276564 160060 276616
rect 276112 276564 276164 276616
rect 117228 276496 117280 276548
rect 226984 276496 227036 276548
rect 51724 275408 51776 275460
rect 182180 275408 182232 275460
rect 57244 275340 57296 275392
rect 187792 275340 187844 275392
rect 61384 275272 61436 275324
rect 194784 275272 194836 275324
rect 124128 271124 124180 271176
rect 208492 271124 208544 271176
rect 161388 265616 161440 265668
rect 252008 265616 252060 265668
rect 245016 259360 245068 259412
rect 580172 259360 580224 259412
rect 3424 255212 3476 255264
rect 68284 255212 68336 255264
rect 119988 254532 120040 254584
rect 222844 254532 222896 254584
rect 582932 245599 582984 245608
rect 582932 245565 582941 245599
rect 582941 245565 582975 245599
rect 582975 245565 582984 245599
rect 582932 245556 582984 245565
rect 133788 243516 133840 243568
rect 258080 243516 258132 243568
rect 258816 243516 258868 243568
rect 329840 243516 329892 243568
rect 3424 241408 3476 241460
rect 53196 241408 53248 241460
rect 147588 238008 147640 238060
rect 268016 238008 268068 238060
rect 233976 219376 234028 219428
rect 579988 219376 580040 219428
rect 3424 188980 3476 189032
rect 65524 188980 65576 189032
rect 231216 179324 231268 179376
rect 580172 179324 580224 179376
rect 3240 164160 3292 164212
rect 148324 164160 148376 164212
rect 233976 163548 234028 163600
rect 316040 163548 316092 163600
rect 148968 163480 149020 163532
rect 269212 163480 269264 163532
rect 3424 150356 3476 150408
rect 71044 150356 71096 150408
rect 3240 137912 3292 137964
rect 21364 137912 21416 137964
rect 582472 126055 582524 126064
rect 582472 126021 582481 126055
rect 582481 126021 582515 126055
rect 582515 126021 582524 126055
rect 582472 126012 582524 126021
rect 162400 113092 162452 113144
rect 580172 113092 580224 113144
rect 3424 111732 3476 111784
rect 141424 111732 141476 111784
rect 3424 97928 3476 97980
rect 53104 97928 53156 97980
rect 350448 93100 350500 93152
rect 414112 93100 414164 93152
rect 472716 91740 472768 91792
rect 490012 91740 490064 91792
rect 3148 85484 3200 85536
rect 3424 71680 3476 71732
rect 142068 71000 142120 71052
rect 263784 71000 263836 71052
rect 162492 60664 162544 60716
rect 579896 60664 579948 60716
rect 3056 59304 3108 59356
rect 3424 45500 3476 45552
rect 255964 36524 256016 36576
rect 303804 36524 303856 36576
rect 162584 33056 162636 33108
rect 580172 33056 580224 33108
rect 162676 20612 162728 20664
rect 580172 20612 580224 20664
rect 129648 17212 129700 17264
rect 255320 17212 255372 17264
rect 126888 13064 126940 13116
rect 252744 13064 252796 13116
rect 245016 12112 245068 12164
rect 306380 12112 306432 12164
rect 228640 12044 228692 12096
rect 324320 12044 324372 12096
rect 230940 11976 230992 12028
rect 327172 11976 327224 12028
rect 224224 11908 224276 11960
rect 321744 11908 321796 11960
rect 223488 11840 223540 11892
rect 323032 11840 323084 11892
rect 342076 11840 342128 11892
rect 158628 11772 158680 11824
rect 276020 11772 276072 11824
rect 144736 11704 144788 11756
rect 266360 11704 266412 11756
rect 342168 11636 342220 11688
rect 169668 10956 169720 11008
rect 244924 10956 244976 11008
rect 165528 10888 165580 10940
rect 251916 10888 251968 10940
rect 179052 10820 179104 10872
rect 291200 10820 291252 10872
rect 176568 10752 176620 10804
rect 288532 10752 288584 10804
rect 136456 10684 136508 10736
rect 249064 10684 249116 10736
rect 154212 10616 154264 10668
rect 273260 10616 273312 10668
rect 140688 10548 140740 10600
rect 263600 10548 263652 10600
rect 128176 10480 128228 10532
rect 251824 10480 251876 10532
rect 252008 10480 252060 10532
rect 309232 10480 309284 10532
rect 85488 10412 85540 10464
rect 223580 10412 223632 10464
rect 268384 10412 268436 10464
rect 353300 10412 353352 10464
rect 162768 10344 162820 10396
rect 580264 10344 580316 10396
rect 3424 10276 3476 10328
rect 149520 9596 149572 9648
rect 269120 9596 269172 9648
rect 153016 9528 153068 9580
rect 271972 9528 272024 9580
rect 145932 9460 145984 9512
rect 267740 9460 267792 9512
rect 142436 9392 142488 9444
rect 265072 9392 265124 9444
rect 138848 9324 138900 9376
rect 262220 9324 262272 9376
rect 122288 9256 122340 9308
rect 249892 9256 249944 9308
rect 118792 9188 118844 9240
rect 247132 9188 247184 9240
rect 267832 9188 267884 9240
rect 335360 9188 335412 9240
rect 115296 9120 115348 9172
rect 245752 9120 245804 9172
rect 269120 9120 269172 9172
rect 345112 9120 345164 9172
rect 108120 9052 108172 9104
rect 240140 9052 240192 9104
rect 258080 9052 258132 9104
rect 342260 9052 342312 9104
rect 111616 8984 111668 9036
rect 242900 8984 242952 9036
rect 264152 8984 264204 9036
rect 352012 8984 352064 9036
rect 104532 8916 104584 8968
rect 237380 8916 237432 8968
rect 240140 8916 240192 8968
rect 334072 8916 334124 8968
rect 156604 8848 156656 8900
rect 274916 8848 274968 8900
rect 160100 8780 160152 8832
rect 277400 8780 277452 8832
rect 171968 8712 172020 8764
rect 233884 8712 233936 8764
rect 233976 8712 234028 8764
rect 327080 8712 327132 8764
rect 237380 8644 237432 8696
rect 320180 8644 320232 8696
rect 177856 8236 177908 8288
rect 289912 8236 289964 8288
rect 167184 8168 167236 8220
rect 283012 8168 283064 8220
rect 170772 8100 170824 8152
rect 285772 8100 285824 8152
rect 163688 8032 163740 8084
rect 280160 8032 280212 8084
rect 135260 7964 135312 8016
rect 259552 7964 259604 8016
rect 131764 7896 131816 7948
rect 256976 7896 257028 7948
rect 77392 7828 77444 7880
rect 218152 7828 218204 7880
rect 73804 7760 73856 7812
rect 215300 7760 215352 7812
rect 343364 7760 343416 7812
rect 409972 7760 410024 7812
rect 38384 7692 38436 7744
rect 180064 7692 180116 7744
rect 181444 7692 181496 7744
rect 292764 7692 292816 7744
rect 304356 7692 304408 7744
rect 380992 7692 381044 7744
rect 70308 7624 70360 7676
rect 212724 7624 212776 7676
rect 298376 7624 298428 7676
rect 376852 7624 376904 7676
rect 66720 7556 66772 7608
rect 209872 7556 209924 7608
rect 292488 7556 292540 7608
rect 371240 7556 371292 7608
rect 377680 7556 377732 7608
rect 434812 7556 434864 7608
rect 174268 7488 174320 7540
rect 287152 7488 287204 7540
rect 184940 7420 184992 7472
rect 295340 7420 295392 7472
rect 188528 7352 188580 7404
rect 298100 7352 298152 7404
rect 192024 7284 192076 7336
rect 300860 7284 300912 7336
rect 195612 7216 195664 7268
rect 303620 7216 303672 7268
rect 199108 7148 199160 7200
rect 305092 7148 305144 7200
rect 202696 7080 202748 7132
rect 307852 7080 307904 7132
rect 206192 7012 206244 7064
rect 310612 7012 310664 7064
rect 63224 6808 63276 6860
rect 207112 6808 207164 6860
rect 215668 6808 215720 6860
rect 317420 6808 317472 6860
rect 59636 6740 59688 6792
rect 205640 6740 205692 6792
rect 212172 6740 212224 6792
rect 314660 6740 314712 6792
rect 56048 6672 56100 6724
rect 202972 6672 203024 6724
rect 208584 6672 208636 6724
rect 311900 6672 311952 6724
rect 52552 6604 52604 6656
rect 200212 6604 200264 6656
rect 205088 6604 205140 6656
rect 309140 6604 309192 6656
rect 48964 6536 49016 6588
rect 197360 6536 197412 6588
rect 201500 6536 201552 6588
rect 307760 6536 307812 6588
rect 44272 6468 44324 6520
rect 194600 6468 194652 6520
rect 197912 6468 197964 6520
rect 305000 6468 305052 6520
rect 40776 6400 40828 6452
rect 191840 6400 191892 6452
rect 194416 6400 194468 6452
rect 302240 6400 302292 6452
rect 345756 6400 345808 6452
rect 411260 6400 411312 6452
rect 37188 6332 37240 6384
rect 189172 6332 189224 6384
rect 190828 6332 190880 6384
rect 299572 6332 299624 6384
rect 339868 6332 339920 6384
rect 407212 6332 407264 6384
rect 33600 6264 33652 6316
rect 186320 6264 186372 6316
rect 187332 6264 187384 6316
rect 296720 6264 296772 6316
rect 335084 6264 335136 6316
rect 403072 6264 403124 6316
rect 8760 6196 8812 6248
rect 168380 6196 168432 6248
rect 173164 6196 173216 6248
rect 287060 6196 287112 6248
rect 318524 6196 318576 6248
rect 392032 6196 392084 6248
rect 4068 6128 4120 6180
rect 165712 6128 165764 6180
rect 169576 6128 169628 6180
rect 284300 6128 284352 6180
rect 307944 6128 307996 6180
rect 383016 6128 383068 6180
rect 445760 6128 445812 6180
rect 483112 6128 483164 6180
rect 101036 6060 101088 6112
rect 234804 6060 234856 6112
rect 271236 6060 271288 6112
rect 357532 6060 357584 6112
rect 126980 5992 127032 6044
rect 254032 5992 254084 6044
rect 274824 5992 274876 6044
rect 360200 5992 360252 6044
rect 130568 5924 130620 5976
rect 256700 5924 256752 5976
rect 278320 5924 278372 5976
rect 362960 5924 363012 5976
rect 162492 5856 162544 5908
rect 278872 5856 278924 5908
rect 166080 5788 166132 5840
rect 281724 5788 281776 5840
rect 176660 5720 176712 5772
rect 289820 5720 289872 5772
rect 180248 5652 180300 5704
rect 292580 5652 292632 5704
rect 183744 5584 183796 5636
rect 293960 5584 294012 5636
rect 69112 5448 69164 5500
rect 212540 5448 212592 5500
rect 303160 5448 303212 5500
rect 380900 5448 380952 5500
rect 65524 5380 65576 5432
rect 209780 5380 209832 5432
rect 292580 5380 292632 5432
rect 372804 5380 372856 5432
rect 62028 5312 62080 5364
rect 207020 5312 207072 5364
rect 288992 5312 289044 5364
rect 369952 5312 370004 5364
rect 58440 5244 58492 5296
rect 204260 5244 204312 5296
rect 285404 5244 285456 5296
rect 367192 5244 367244 5296
rect 54944 5176 54996 5228
rect 201592 5176 201644 5228
rect 216864 5176 216916 5228
rect 276664 5176 276716 5228
rect 281908 5176 281960 5228
rect 365720 5176 365772 5228
rect 51356 5108 51408 5160
rect 199016 5108 199068 5160
rect 209780 5108 209832 5160
rect 295984 5108 296036 5160
rect 296076 5108 296128 5160
rect 375380 5108 375432 5160
rect 26516 5040 26568 5092
rect 180892 5040 180944 5092
rect 257068 5040 257120 5092
rect 347780 5040 347832 5092
rect 30104 4972 30156 5024
rect 183652 4972 183704 5024
rect 260656 4972 260708 5024
rect 350540 4972 350592 5024
rect 21824 4904 21876 4956
rect 178040 4904 178092 4956
rect 253480 4904 253532 4956
rect 345020 4904 345072 4956
rect 17040 4836 17092 4888
rect 173992 4836 174044 4888
rect 246396 4836 246448 4888
rect 339592 4836 339644 4888
rect 384764 4836 384816 4888
rect 438952 4836 439004 4888
rect 12348 4768 12400 4820
rect 171140 4768 171192 4820
rect 242900 4768 242952 4820
rect 337016 4768 337068 4820
rect 370596 4768 370648 4820
rect 429200 4768 429252 4820
rect 72608 4700 72660 4752
rect 214012 4700 214064 4752
rect 299664 4700 299716 4752
rect 378140 4700 378192 4752
rect 79692 4632 79744 4684
rect 219532 4632 219584 4684
rect 306748 4632 306800 4684
rect 383752 4632 383804 4684
rect 76196 4564 76248 4616
rect 216956 4564 217008 4616
rect 310244 4564 310296 4616
rect 385132 4564 385184 4616
rect 86868 4496 86920 4548
rect 224960 4496 225012 4548
rect 317328 4496 317380 4548
rect 390744 4496 390796 4548
rect 83280 4428 83332 4480
rect 222200 4428 222252 4480
rect 313832 4428 313884 4480
rect 387892 4428 387944 4480
rect 90364 4360 90416 4412
rect 227720 4360 227772 4412
rect 320916 4360 320968 4412
rect 393320 4360 393372 4412
rect 93952 4292 94004 4344
rect 229192 4292 229244 4344
rect 328000 4292 328052 4344
rect 398840 4292 398892 4344
rect 97448 4224 97500 4276
rect 231952 4224 232004 4276
rect 324412 4224 324464 4276
rect 396080 4224 396132 4276
rect 14740 4088 14792 4140
rect 18604 4088 18656 4140
rect 18236 4020 18288 4072
rect 33784 4088 33836 4140
rect 25320 4020 25372 4072
rect 29644 4020 29696 4072
rect 32404 4020 32456 4072
rect 36544 4088 36596 4140
rect 34796 4020 34848 4072
rect 57244 4088 57296 4140
rect 67916 4088 67968 4140
rect 195244 4088 195296 4140
rect 214472 4088 214524 4140
rect 229836 4088 229888 4140
rect 233976 4088 234028 4140
rect 237012 4088 237064 4140
rect 54484 4020 54536 4072
rect 60832 4020 60884 4072
rect 192484 4020 192536 4072
rect 207388 4020 207440 4072
rect 313924 4088 313976 4140
rect 316224 4088 316276 4140
rect 389824 4088 389876 4140
rect 393044 4088 393096 4140
rect 393964 4088 394016 4140
rect 400220 4088 400272 4140
rect 401324 4088 401376 4140
rect 402520 4088 402572 4140
rect 402980 4088 403032 4140
rect 451280 4088 451332 4140
rect 456892 4088 456944 4140
rect 461584 4088 461636 4140
rect 474004 4088 474056 4140
rect 497096 4088 497148 4140
rect 501604 4088 501656 4140
rect 556160 4088 556212 4140
rect 558276 4088 558328 4140
rect 240784 4020 240836 4072
rect 247592 4020 247644 4072
rect 273904 4020 273956 4072
rect 280712 4020 280764 4072
rect 287796 4020 287848 4072
rect 1676 3952 1728 4004
rect 22744 3952 22796 4004
rect 27712 3952 27764 4004
rect 51724 3952 51776 4004
rect 53748 3952 53800 4004
rect 191104 3952 191156 4004
rect 210976 3952 211028 4004
rect 250444 3952 250496 4004
rect 258172 3952 258224 4004
rect 258816 3952 258868 4004
rect 265348 3952 265400 4004
rect 268384 3952 268436 4004
rect 272432 3952 272484 4004
rect 282184 3952 282236 4004
rect 283104 3952 283156 4004
rect 291292 3952 291344 4004
rect 291384 3952 291436 4004
rect 293224 3952 293276 4004
rect 294880 4020 294932 4072
rect 374000 4020 374052 4072
rect 383568 4020 383620 4072
rect 384304 4020 384356 4072
rect 385960 4020 386012 4072
rect 388444 4020 388496 4072
rect 389456 4020 389508 4072
rect 369860 3952 369912 4004
rect 382372 3952 382424 4004
rect 437664 3952 437716 4004
rect 13544 3884 13596 3936
rect 39304 3884 39356 3936
rect 43076 3884 43128 3936
rect 193220 3884 193272 3936
rect 218060 3884 218112 3936
rect 262864 3884 262916 3936
rect 266544 3884 266596 3936
rect 349804 3884 349856 3936
rect 352840 3884 352892 3936
rect 353944 3884 353996 3936
rect 356336 3884 356388 3936
rect 357348 3884 357400 3936
rect 357532 3884 357584 3936
rect 358728 3884 358780 3936
rect 7656 3816 7708 3868
rect 32312 3816 32364 3868
rect 35992 3816 36044 3868
rect 187700 3816 187752 3868
rect 203892 3816 203944 3868
rect 252008 3816 252060 3868
rect 254676 3816 254728 3868
rect 2872 3748 2924 3800
rect 25504 3748 25556 3800
rect 28908 3748 28960 3800
rect 183560 3748 183612 3800
rect 196808 3748 196860 3800
rect 255964 3748 256016 3800
rect 261760 3816 261812 3868
rect 278044 3816 278096 3868
rect 279516 3816 279568 3868
rect 286324 3816 286376 3868
rect 269120 3748 269172 3800
rect 273628 3748 273680 3800
rect 355232 3748 355284 3800
rect 356704 3748 356756 3800
rect 358636 3816 358688 3868
rect 420920 3884 420972 3936
rect 424324 3884 424376 3936
rect 431224 3884 431276 3936
rect 375196 3816 375248 3868
rect 431960 3816 432012 3868
rect 446220 4020 446272 4072
rect 460204 4020 460256 4072
rect 462780 4020 462832 4072
rect 486332 4020 486384 4072
rect 440332 3952 440384 4004
rect 459192 3952 459244 4004
rect 485044 3952 485096 4004
rect 563244 3952 563296 4004
rect 568580 3952 568632 4004
rect 467104 3884 467156 3936
rect 468668 3884 468720 3936
rect 476764 3884 476816 3936
rect 479340 3884 479392 3936
rect 480904 3884 480956 3936
rect 508504 3884 508556 3936
rect 443092 3816 443144 3868
rect 447140 3816 447192 3868
rect 469864 3816 469916 3868
rect 504180 3816 504232 3868
rect 512644 3816 512696 3868
rect 363604 3748 363656 3800
rect 368204 3748 368256 3800
rect 427912 3748 427964 3800
rect 468484 3748 468536 3800
rect 493508 3748 493560 3800
rect 504364 3748 504416 3800
rect 19432 3680 19484 3732
rect 176752 3680 176804 3732
rect 189724 3680 189776 3732
rect 253204 3680 253256 3732
rect 259460 3680 259512 3732
rect 349160 3680 349212 3732
rect 354036 3680 354088 3732
rect 416780 3680 416832 3732
rect 420184 3680 420236 3732
rect 421380 3680 421432 3732
rect 464436 3680 464488 3732
rect 473452 3680 473504 3732
rect 493416 3680 493468 3732
rect 498200 3680 498252 3732
rect 503720 3680 503772 3732
rect 539600 3680 539652 3732
rect 550916 3680 550968 3732
rect 572 3612 624 3664
rect 14464 3612 14516 3664
rect 20628 3612 20680 3664
rect 176936 3612 176988 3664
rect 200304 3612 200356 3664
rect 246304 3612 246356 3664
rect 248788 3612 248840 3664
rect 249708 3612 249760 3664
rect 252376 3612 252428 3664
rect 342904 3612 342956 3664
rect 351644 3612 351696 3664
rect 415400 3612 415452 3664
rect 421564 3612 421616 3664
rect 424968 3612 425020 3664
rect 467840 3612 467892 3664
rect 475384 3612 475436 3664
rect 476948 3612 477000 3664
rect 502892 3612 502944 3664
rect 11152 3544 11204 3596
rect 169760 3544 169812 3596
rect 182548 3544 182600 3596
rect 209044 3544 209096 3596
rect 213368 3544 213420 3596
rect 215944 3544 215996 3596
rect 221556 3544 221608 3596
rect 224224 3544 224276 3596
rect 225144 3544 225196 3596
rect 228640 3544 228692 3596
rect 228732 3544 228784 3596
rect 230940 3544 230992 3596
rect 231032 3544 231084 3596
rect 322020 3544 322072 3596
rect 322112 3544 322164 3596
rect 324964 3544 325016 3596
rect 394700 3544 394752 3596
rect 395344 3544 395396 3596
rect 396724 3544 396776 3596
rect 397736 3544 397788 3596
rect 399484 3544 399536 3596
rect 443828 3544 443880 3596
rect 444288 3544 444340 3596
rect 448612 3544 448664 3596
rect 450544 3544 450596 3596
rect 472624 3544 472676 3596
rect 474556 3544 474608 3596
rect 9956 3476 10008 3528
rect 164884 3476 164936 3528
rect 165528 3476 165580 3528
rect 168380 3476 168432 3528
rect 169668 3476 169720 3528
rect 175464 3476 175516 3528
rect 176568 3476 176620 3528
rect 193220 3476 193272 3528
rect 5264 3408 5316 3460
rect 165804 3408 165856 3460
rect 186136 3408 186188 3460
rect 222752 3476 222804 3528
rect 223488 3476 223540 3528
rect 223948 3476 224000 3528
rect 224868 3476 224920 3528
rect 234068 3476 234120 3528
rect 234620 3476 234672 3528
rect 239312 3476 239364 3528
rect 240140 3476 240192 3528
rect 241704 3476 241756 3528
rect 242808 3476 242860 3528
rect 245200 3476 245252 3528
rect 338304 3476 338356 3528
rect 338672 3476 338724 3528
rect 339408 3476 339460 3528
rect 340972 3476 341024 3528
rect 341984 3476 342036 3528
rect 348056 3476 348108 3528
rect 349068 3476 349120 3528
rect 349252 3476 349304 3528
rect 350448 3476 350500 3528
rect 404820 3476 404872 3528
rect 405648 3476 405700 3528
rect 406016 3476 406068 3528
rect 407028 3476 407080 3528
rect 407212 3476 407264 3528
rect 409144 3476 409196 3528
rect 409604 3476 409656 3528
rect 410524 3476 410576 3528
rect 411904 3476 411956 3528
rect 412548 3476 412600 3528
rect 413100 3476 413152 3528
rect 413928 3476 413980 3528
rect 414296 3476 414348 3528
rect 415308 3476 415360 3528
rect 416688 3476 416740 3528
rect 417424 3476 417476 3528
rect 418988 3476 419040 3528
rect 419448 3476 419500 3528
rect 461032 3476 461084 3528
rect 471060 3476 471112 3528
rect 471888 3476 471940 3528
rect 478144 3476 478196 3528
rect 479524 3476 479576 3528
rect 481732 3544 481784 3596
rect 482928 3544 482980 3596
rect 485228 3544 485280 3596
rect 485688 3544 485740 3596
rect 486424 3544 486476 3596
rect 487068 3544 487120 3596
rect 487620 3544 487672 3596
rect 489184 3544 489236 3596
rect 510620 3612 510672 3664
rect 505376 3544 505428 3596
rect 519544 3612 519596 3664
rect 518348 3544 518400 3596
rect 535552 3612 535604 3664
rect 554964 3612 555016 3664
rect 558184 3612 558236 3664
rect 566832 3612 566884 3664
rect 570144 3612 570196 3664
rect 533712 3544 533764 3596
rect 546592 3544 546644 3596
rect 546684 3544 546736 3596
rect 548524 3544 548576 3596
rect 551468 3544 551520 3596
rect 556804 3544 556856 3596
rect 559748 3544 559800 3596
rect 566004 3544 566056 3596
rect 570328 3544 570380 3596
rect 572720 3544 572772 3596
rect 501788 3476 501840 3528
rect 502248 3476 502300 3528
rect 502984 3476 503036 3528
rect 503628 3476 503680 3528
rect 507676 3476 507728 3528
rect 528652 3476 528704 3528
rect 529020 3476 529072 3528
rect 529848 3476 529900 3528
rect 532516 3476 532568 3528
rect 533344 3476 533396 3528
rect 534908 3476 534960 3528
rect 535368 3476 535420 3528
rect 536104 3476 536156 3528
rect 536748 3476 536800 3528
rect 537208 3476 537260 3528
rect 538128 3476 538180 3528
rect 538404 3476 538456 3528
rect 539508 3476 539560 3528
rect 541992 3476 542044 3528
rect 543004 3476 543056 3528
rect 543188 3476 543240 3528
rect 544292 3476 544344 3528
rect 544384 3476 544436 3528
rect 545028 3476 545080 3528
rect 545488 3476 545540 3528
rect 547144 3476 547196 3528
rect 550272 3476 550324 3528
rect 551284 3476 551336 3528
rect 553768 3476 553820 3528
rect 554688 3476 554740 3528
rect 560852 3476 560904 3528
rect 561588 3476 561640 3528
rect 562048 3476 562100 3528
rect 562968 3476 563020 3528
rect 564440 3476 564492 3528
rect 566464 3476 566516 3528
rect 568028 3476 568080 3528
rect 569224 3476 569276 3528
rect 571524 3476 571576 3528
rect 572628 3476 572680 3528
rect 577412 3476 577464 3528
rect 578240 3476 578292 3528
rect 583392 3476 583444 3528
rect 23020 3340 23072 3392
rect 6460 3272 6512 3324
rect 7564 3272 7616 3324
rect 24216 3272 24268 3324
rect 31300 3272 31352 3324
rect 41880 3340 41932 3392
rect 58624 3340 58676 3392
rect 75000 3340 75052 3392
rect 196624 3340 196676 3392
rect 219256 3340 219308 3392
rect 39580 3272 39632 3324
rect 43444 3272 43496 3324
rect 45468 3272 45520 3324
rect 61384 3272 61436 3324
rect 80888 3272 80940 3324
rect 81348 3272 81400 3324
rect 84476 3272 84528 3324
rect 85488 3272 85540 3324
rect 87604 3272 87656 3324
rect 87972 3272 88024 3324
rect 88984 3272 89036 3324
rect 35164 3204 35216 3256
rect 40684 3204 40736 3256
rect 82084 3204 82136 3256
rect 199384 3272 199436 3324
rect 91560 3204 91612 3256
rect 93124 3204 93176 3256
rect 15936 3136 15988 3188
rect 17224 3136 17276 3188
rect 50160 3136 50212 3188
rect 86224 3136 86276 3188
rect 57244 3068 57296 3120
rect 85672 3068 85724 3120
rect 200764 3204 200816 3256
rect 238024 3408 238076 3460
rect 238116 3408 238168 3460
rect 326804 3408 326856 3460
rect 329104 3408 329156 3460
rect 331588 3408 331640 3460
rect 332508 3408 332560 3460
rect 337476 3408 337528 3460
rect 405832 3408 405884 3460
rect 408408 3408 408460 3460
rect 231124 3340 231176 3392
rect 226340 3272 226392 3324
rect 227628 3272 227680 3324
rect 93308 3068 93360 3120
rect 203524 3136 203576 3188
rect 237380 3340 237432 3392
rect 240508 3340 240560 3392
rect 267832 3340 267884 3392
rect 270040 3340 270092 3392
rect 298468 3340 298520 3392
rect 299388 3340 299440 3392
rect 305552 3340 305604 3392
rect 306288 3340 306340 3392
rect 312636 3340 312688 3392
rect 313188 3340 313240 3392
rect 323308 3340 323360 3392
rect 329196 3340 329248 3392
rect 331864 3340 331916 3392
rect 350448 3340 350500 3392
rect 352564 3340 352616 3392
rect 358820 3340 358872 3392
rect 363512 3340 363564 3392
rect 364248 3340 364300 3392
rect 364616 3340 364668 3392
rect 366364 3340 366416 3392
rect 367008 3340 367060 3392
rect 367744 3340 367796 3392
rect 371700 3340 371752 3392
rect 373264 3340 373316 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 376484 3340 376536 3392
rect 377404 3340 377456 3392
rect 378876 3340 378928 3392
rect 379428 3340 379480 3392
rect 381176 3340 381228 3392
rect 382924 3340 382976 3392
rect 423772 3340 423824 3392
rect 425796 3340 425848 3392
rect 427268 3340 427320 3392
rect 428464 3340 428516 3392
rect 429660 3340 429712 3392
rect 430488 3340 430540 3392
rect 430856 3340 430908 3392
rect 431868 3340 431920 3392
rect 432052 3340 432104 3392
rect 433248 3340 433300 3392
rect 233424 3272 233476 3324
rect 258172 3272 258224 3324
rect 258264 3272 258316 3324
rect 260104 3272 260156 3324
rect 277124 3272 277176 3324
rect 307024 3272 307076 3324
rect 309048 3272 309100 3324
rect 385040 3272 385092 3324
rect 388260 3272 388312 3324
rect 389916 3272 389968 3324
rect 390652 3272 390704 3324
rect 391756 3272 391808 3324
rect 391848 3272 391900 3324
rect 392584 3272 392636 3324
rect 436652 3340 436704 3392
rect 436744 3340 436796 3392
rect 437388 3340 437440 3392
rect 439136 3340 439188 3392
rect 440148 3340 440200 3392
rect 456064 3408 456116 3460
rect 460388 3408 460440 3460
rect 462964 3408 463016 3460
rect 463976 3408 464028 3460
rect 452108 3340 452160 3392
rect 453304 3340 453356 3392
rect 434444 3272 434496 3324
rect 435364 3272 435416 3324
rect 437940 3272 437992 3324
rect 440884 3272 440936 3324
rect 441528 3272 441580 3324
rect 446404 3272 446456 3324
rect 447416 3272 447468 3324
rect 456984 3340 457036 3392
rect 461584 3340 461636 3392
rect 455696 3272 455748 3324
rect 472716 3340 472768 3392
rect 480536 3340 480588 3392
rect 482284 3340 482336 3392
rect 488816 3340 488868 3392
rect 489828 3340 489880 3392
rect 492312 3408 492364 3460
rect 493324 3408 493376 3460
rect 494704 3408 494756 3460
rect 495348 3408 495400 3460
rect 495900 3408 495952 3460
rect 496728 3408 496780 3460
rect 499396 3408 499448 3460
rect 497004 3340 497056 3392
rect 511264 3408 511316 3460
rect 511908 3408 511960 3460
rect 512460 3408 512512 3460
rect 513288 3408 513340 3460
rect 513564 3408 513616 3460
rect 514668 3408 514720 3460
rect 514760 3408 514812 3460
rect 515864 3408 515916 3460
rect 519544 3408 519596 3460
rect 520188 3408 520240 3460
rect 520740 3408 520792 3460
rect 521568 3408 521620 3460
rect 521844 3408 521896 3460
rect 522948 3408 523000 3460
rect 524236 3408 524288 3460
rect 525156 3408 525208 3460
rect 526628 3408 526680 3460
rect 527088 3408 527140 3460
rect 527824 3408 527876 3460
rect 542360 3408 542412 3460
rect 552664 3408 552716 3460
rect 560392 3408 560444 3460
rect 576308 3408 576360 3460
rect 576768 3408 576820 3460
rect 521936 3340 521988 3392
rect 523040 3340 523092 3392
rect 525064 3340 525116 3392
rect 531320 3340 531372 3392
rect 533436 3340 533488 3392
rect 472256 3272 472308 3324
rect 478052 3272 478104 3324
rect 482836 3272 482888 3324
rect 510068 3272 510120 3324
rect 518164 3272 518216 3324
rect 235816 3204 235868 3256
rect 232228 3136 232280 3188
rect 233148 3136 233200 3188
rect 245016 3204 245068 3256
rect 255872 3204 255924 3256
rect 323584 3204 323636 3256
rect 330392 3204 330444 3256
rect 398932 3204 398984 3256
rect 400864 3204 400916 3256
rect 403624 3204 403676 3256
rect 452660 3204 452712 3256
rect 453304 3204 453356 3256
rect 460296 3204 460348 3256
rect 506480 3204 506532 3256
rect 507768 3204 507820 3256
rect 242164 3136 242216 3188
rect 249984 3136 250036 3188
rect 258080 3136 258132 3188
rect 262956 3136 263008 3188
rect 320824 3136 320876 3188
rect 325608 3136 325660 3188
rect 340144 3136 340196 3188
rect 344560 3136 344612 3188
rect 407764 3136 407816 3188
rect 410800 3136 410852 3188
rect 454776 3136 454828 3188
rect 465172 3136 465224 3188
rect 466368 3136 466420 3188
rect 469864 3136 469916 3188
rect 471244 3136 471296 3188
rect 530124 3136 530176 3188
rect 531228 3136 531280 3188
rect 569132 3136 569184 3188
rect 572904 3136 572956 3188
rect 98644 3068 98696 3120
rect 99288 3068 99340 3120
rect 102232 3068 102284 3120
rect 105544 3068 105596 3120
rect 105728 3068 105780 3120
rect 106188 3068 106240 3120
rect 110512 3068 110564 3120
rect 111708 3068 111760 3120
rect 112812 3068 112864 3120
rect 115112 3068 115164 3120
rect 116400 3068 116452 3120
rect 117228 3068 117280 3120
rect 117596 3068 117648 3120
rect 118608 3068 118660 3120
rect 214564 3068 214616 3120
rect 244096 3068 244148 3120
rect 267004 3068 267056 3120
rect 268844 3068 268896 3120
rect 280804 3068 280856 3120
rect 284300 3068 284352 3120
rect 300124 3068 300176 3120
rect 71504 3000 71556 3052
rect 106924 3000 106976 3052
rect 109316 3000 109368 3052
rect 112444 3000 112496 3052
rect 114008 3000 114060 3052
rect 221464 3000 221516 3052
rect 251180 3000 251232 3052
rect 258724 3000 258776 3052
rect 276020 3000 276072 3052
rect 284944 3000 284996 3052
rect 286600 3000 286652 3052
rect 289084 3000 289136 3052
rect 290188 3000 290240 3052
rect 292488 3000 292540 3052
rect 293684 3000 293736 3052
rect 311440 3068 311492 3120
rect 64328 2932 64380 2984
rect 46664 2864 46716 2916
rect 50344 2864 50396 2916
rect 78588 2864 78640 2916
rect 89168 2932 89220 2984
rect 97264 2932 97316 2984
rect 99840 2932 99892 2984
rect 206284 2932 206336 2984
rect 267740 2932 267792 2984
rect 271144 2932 271196 2984
rect 297272 2932 297324 2984
rect 298376 2932 298428 2984
rect 300768 2932 300820 2984
rect 314016 3000 314068 3052
rect 315028 3000 315080 3052
rect 318064 3000 318116 3052
rect 334164 3068 334216 3120
rect 361120 3068 361172 3120
rect 336004 3000 336056 3052
rect 336280 3000 336332 3052
rect 360844 3000 360896 3052
rect 362316 3000 362368 3052
rect 364984 3000 365036 3052
rect 365812 3000 365864 3052
rect 415492 3068 415544 3120
rect 422576 3068 422628 3120
rect 464344 3068 464396 3120
rect 573916 3068 573968 3120
rect 575572 3068 575624 3120
rect 420092 3000 420144 3052
rect 428464 3000 428516 3052
rect 316684 2932 316736 2984
rect 332692 2932 332744 2984
rect 346860 2932 346912 2984
rect 346952 2932 347004 2984
rect 372896 2932 372948 2984
rect 425704 2932 425756 2984
rect 426164 2932 426216 2984
rect 433248 2932 433300 2984
rect 435548 2932 435600 2984
rect 90272 2864 90324 2916
rect 92756 2864 92808 2916
rect 93308 2864 93360 2916
rect 96252 2864 96304 2916
rect 101404 2864 101456 2916
rect 103336 2864 103388 2916
rect 94504 2796 94556 2848
rect 106924 2864 106976 2916
rect 108304 2796 108356 2848
rect 121092 2796 121144 2848
rect 221648 2864 221700 2916
rect 301964 2864 302016 2916
rect 379704 2864 379756 2916
rect 379980 2864 380032 2916
rect 387156 2864 387208 2916
rect 394240 2864 394292 2916
rect 442264 2864 442316 2916
rect 442632 3000 442684 3052
rect 447784 3000 447836 3052
rect 454500 3000 454552 3052
rect 475752 3000 475804 3052
rect 479616 3000 479668 3052
rect 547880 3000 547932 3052
rect 555424 3000 555476 3052
rect 558552 3000 558604 3052
rect 564624 3000 564676 3052
rect 578608 3000 578660 3052
rect 579620 3000 579672 3052
rect 445024 2932 445076 2984
rect 445760 2932 445812 2984
rect 489920 2932 489972 2984
rect 497464 2932 497516 2984
rect 525432 2932 525484 2984
rect 526444 2932 526496 2984
rect 572720 2932 572772 2984
rect 574192 2932 574244 2984
rect 449164 2864 449216 2916
rect 123484 2796 123536 2848
rect 124128 2796 124180 2848
rect 124680 2796 124732 2848
rect 125416 2796 125468 2848
rect 125876 2796 125928 2848
rect 126888 2796 126940 2848
rect 132960 2796 133012 2848
rect 133788 2796 133840 2848
rect 134156 2796 134208 2848
rect 135168 2796 135220 2848
rect 140044 2796 140096 2848
rect 140688 2796 140740 2848
rect 141240 2796 141292 2848
rect 142068 2796 142120 2848
rect 143540 2796 143592 2848
rect 144828 2796 144880 2848
rect 147128 2796 147180 2848
rect 147588 2796 147640 2848
rect 148324 2796 148376 2848
rect 148968 2796 149020 2848
rect 150624 2796 150676 2848
rect 151728 2796 151780 2848
rect 151820 2796 151872 2848
rect 153108 2796 153160 2848
rect 155408 2796 155460 2848
rect 155868 2796 155920 2848
rect 157800 2796 157852 2848
rect 158628 2796 158680 2848
rect 158904 2796 158956 2848
rect 160008 2796 160060 2848
rect 169852 2796 169904 2848
rect 302884 2796 302936 2848
rect 396540 2796 396592 2848
rect 412732 2796 412784 2848
rect 417884 2796 417936 2848
rect 454684 2796 454736 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 141424 703656 141476 703662
rect 141424 703598 141476 703604
rect 3424 700392 3476 700398
rect 3424 700334 3476 700340
rect 3056 672036 3108 672042
rect 3056 671978 3108 671984
rect 3068 671265 3096 671978
rect 3054 671256 3110 671265
rect 3054 671191 3110 671200
rect 3332 619608 3384 619614
rect 3332 619550 3384 619556
rect 3344 619177 3372 619550
rect 3330 619168 3386 619177
rect 3330 619103 3386 619112
rect 3240 607164 3292 607170
rect 3240 607106 3292 607112
rect 3252 606121 3280 607106
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3240 463684 3292 463690
rect 3240 463626 3292 463632
rect 3252 462641 3280 463626
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3240 398812 3292 398818
rect 3240 398754 3292 398760
rect 3252 397497 3280 398754
rect 3238 397488 3294 397497
rect 3238 397423 3294 397432
rect 3436 358465 3464 700334
rect 8128 699786 8156 703520
rect 14464 702432 14516 702438
rect 14464 702374 14516 702380
rect 8116 699780 8168 699786
rect 8116 699722 8168 699728
rect 3516 658232 3568 658238
rect 3514 658200 3516 658209
rect 3568 658200 3570 658209
rect 3514 658135 3570 658144
rect 3514 633312 3570 633321
rect 3514 633247 3570 633256
rect 3528 632097 3556 633247
rect 3514 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 580952 3570 580961
rect 3514 580887 3570 580896
rect 3528 580009 3556 580887
rect 3514 580000 3570 580009
rect 3514 579935 3570 579944
rect 3516 567180 3568 567186
rect 3516 567122 3568 567128
rect 3528 566953 3556 567122
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3516 554736 3568 554742
rect 3516 554678 3568 554684
rect 3528 553897 3556 554678
rect 3514 553888 3570 553897
rect 3514 553823 3570 553832
rect 3516 516112 3568 516118
rect 3516 516054 3568 516060
rect 3528 514865 3556 516054
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 14476 502314 14504 702374
rect 17224 702364 17276 702370
rect 17224 702306 17276 702312
rect 14556 699712 14608 699718
rect 14556 699654 14608 699660
rect 14568 658238 14596 699654
rect 14556 658232 14608 658238
rect 14556 658174 14608 658180
rect 3516 502308 3568 502314
rect 3516 502250 3568 502256
rect 14464 502308 14516 502314
rect 14464 502250 14516 502256
rect 3528 501809 3556 502250
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 17236 449886 17264 702306
rect 18602 701312 18658 701321
rect 18602 701247 18658 701256
rect 17224 449880 17276 449886
rect 17224 449822 17276 449828
rect 3516 423632 3568 423638
rect 3514 423600 3516 423609
rect 3568 423600 3570 423609
rect 3514 423535 3570 423544
rect 18616 398818 18644 701247
rect 21362 700768 21418 700777
rect 21362 700703 21418 700712
rect 18604 398812 18656 398818
rect 18604 398754 18656 398760
rect 3516 372564 3568 372570
rect 3516 372506 3568 372512
rect 3528 371385 3556 372506
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 3424 306332 3476 306338
rect 3424 306274 3476 306280
rect 3436 306241 3464 306274
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 3068 293185 3096 293898
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 18604 279608 18656 279614
rect 18604 279550 18656 279556
rect 17224 279540 17276 279546
rect 17224 279482 17276 279488
rect 7564 279472 7616 279478
rect 7564 279414 7616 279420
rect 3424 255264 3476 255270
rect 3424 255206 3476 255212
rect 3436 254153 3464 255206
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3424 241460 3476 241466
rect 3424 241402 3476 241408
rect 3436 241097 3464 241402
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3422 202872 3478 202881
rect 3422 202807 3478 202816
rect 3436 201929 3464 202807
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3330 33144 3386 33153
rect 3330 33079 3386 33088
rect 3344 32473 3372 33079
rect 3330 32464 3386 32473
rect 3330 32399 3386 32408
rect 3422 20632 3478 20641
rect 3422 20567 3478 20576
rect 3436 19417 3464 20567
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 10328 3476 10334
rect 3424 10270 3476 10276
rect 3436 6497 3464 10270
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 572 3664 624 3670
rect 572 3606 624 3612
rect 584 480 612 3606
rect 1688 480 1716 3946
rect 2872 3800 2924 3806
rect 2872 3742 2924 3748
rect 2884 480 2912 3742
rect 4080 480 4108 6122
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 7576 3330 7604 279414
rect 14464 278044 14516 278050
rect 14464 277986 14516 277992
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 7656 3868 7708 3874
rect 7656 3810 7708 3816
rect 6460 3324 6512 3330
rect 6460 3266 6512 3272
rect 7564 3324 7616 3330
rect 7564 3266 7616 3272
rect 6472 480 6500 3266
rect 7668 480 7696 3810
rect 8772 480 8800 6190
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9968 480 9996 3470
rect 11164 480 11192 3538
rect 12360 480 12388 4762
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 480 13584 3878
rect 14476 3670 14504 277986
rect 17040 4888 17092 4894
rect 17040 4830 17092 4836
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14464 3664 14516 3670
rect 14464 3606 14516 3612
rect 14752 480 14780 4082
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15948 480 15976 3130
rect 17052 480 17080 4830
rect 17236 3194 17264 279482
rect 18616 4146 18644 279550
rect 21376 137970 21404 700703
rect 24320 699990 24348 703520
rect 29642 701176 29698 701185
rect 29642 701111 29698 701120
rect 24308 699984 24360 699990
rect 24308 699926 24360 699932
rect 29656 306338 29684 701111
rect 40512 701049 40540 703520
rect 71044 702092 71096 702098
rect 71044 702034 71096 702040
rect 65524 702024 65576 702030
rect 65524 701966 65576 701972
rect 40498 701040 40554 701049
rect 40498 700975 40554 700984
rect 53104 700528 53156 700534
rect 53104 700470 53156 700476
rect 32402 700088 32458 700097
rect 32402 700023 32458 700032
rect 35164 700052 35216 700058
rect 32416 463690 32444 700023
rect 35164 699994 35216 700000
rect 35176 672042 35204 699994
rect 40684 699916 40736 699922
rect 40684 699858 40736 699864
rect 35164 672036 35216 672042
rect 35164 671978 35216 671984
rect 40696 607170 40724 699858
rect 43444 699848 43496 699854
rect 43444 699790 43496 699796
rect 40684 607164 40736 607170
rect 40684 607106 40736 607112
rect 43456 554742 43484 699790
rect 43444 554736 43496 554742
rect 43444 554678 43496 554684
rect 32404 463684 32456 463690
rect 32404 463626 32456 463632
rect 29644 306332 29696 306338
rect 29644 306274 29696 306280
rect 35164 279948 35216 279954
rect 35164 279890 35216 279896
rect 29644 279676 29696 279682
rect 29644 279618 29696 279624
rect 25504 278316 25556 278322
rect 25504 278258 25556 278264
rect 22744 278180 22796 278186
rect 22744 278122 22796 278128
rect 21364 137964 21416 137970
rect 21364 137906 21416 137912
rect 21824 4956 21876 4962
rect 21824 4898 21876 4904
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 18248 480 18276 4014
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19444 480 19472 3674
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 20640 480 20668 3606
rect 21836 480 21864 4898
rect 22756 4010 22784 278122
rect 25320 4072 25372 4078
rect 25320 4014 25372 4020
rect 22744 4004 22796 4010
rect 22744 3946 22796 3952
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 23032 480 23060 3334
rect 24216 3324 24268 3330
rect 24216 3266 24268 3272
rect 24228 480 24256 3266
rect 25332 480 25360 4014
rect 25516 3806 25544 278258
rect 26516 5092 26568 5098
rect 26516 5034 26568 5040
rect 25504 3800 25556 3806
rect 25504 3742 25556 3748
rect 26528 480 26556 5034
rect 29656 4078 29684 279618
rect 32404 278520 32456 278526
rect 32404 278462 32456 278468
rect 32416 6914 32444 278462
rect 33784 276684 33836 276690
rect 33784 276626 33836 276632
rect 32324 6886 32444 6914
rect 30104 5024 30156 5030
rect 30104 4966 30156 4972
rect 29644 4072 29696 4078
rect 29644 4014 29696 4020
rect 27712 4004 27764 4010
rect 27712 3946 27764 3952
rect 27724 480 27752 3946
rect 28908 3800 28960 3806
rect 28908 3742 28960 3748
rect 28920 480 28948 3742
rect 30116 480 30144 4966
rect 32324 3874 32352 6886
rect 33600 6316 33652 6322
rect 33600 6258 33652 6264
rect 32404 4072 32456 4078
rect 32404 4014 32456 4020
rect 32312 3868 32364 3874
rect 32312 3810 32364 3816
rect 31300 3324 31352 3330
rect 31300 3266 31352 3272
rect 31312 480 31340 3266
rect 32416 480 32444 4014
rect 33612 480 33640 6258
rect 33796 4146 33824 276626
rect 33784 4140 33836 4146
rect 33784 4082 33836 4088
rect 34796 4072 34848 4078
rect 34796 4014 34848 4020
rect 34808 480 34836 4014
rect 35176 3262 35204 279890
rect 50344 279880 50396 279886
rect 50344 279822 50396 279828
rect 43444 279812 43496 279818
rect 43444 279754 43496 279760
rect 36544 279744 36596 279750
rect 36544 279686 36596 279692
rect 36556 4146 36584 279686
rect 39304 278656 39356 278662
rect 39304 278598 39356 278604
rect 38384 7744 38436 7750
rect 38384 7686 38436 7692
rect 37188 6384 37240 6390
rect 37188 6326 37240 6332
rect 36544 4140 36596 4146
rect 36544 4082 36596 4088
rect 35992 3868 36044 3874
rect 35992 3810 36044 3816
rect 35164 3256 35216 3262
rect 35164 3198 35216 3204
rect 36004 480 36032 3810
rect 37200 480 37228 6326
rect 38396 480 38424 7686
rect 39316 3942 39344 278598
rect 40684 276752 40736 276758
rect 40684 276694 40736 276700
rect 39304 3936 39356 3942
rect 39304 3878 39356 3884
rect 39580 3324 39632 3330
rect 39580 3266 39632 3272
rect 39592 480 39620 3266
rect 40696 3262 40724 276694
rect 40776 6452 40828 6458
rect 40776 6394 40828 6400
rect 40684 3256 40736 3262
rect 40684 3198 40736 3204
rect 40788 3074 40816 6394
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 40696 3046 40816 3074
rect 40696 480 40724 3046
rect 41892 480 41920 3334
rect 43088 480 43116 3878
rect 43456 3330 43484 279754
rect 48228 278112 48280 278118
rect 48228 278054 48280 278060
rect 48240 6914 48268 278054
rect 47872 6886 48268 6914
rect 44272 6520 44324 6526
rect 44272 6462 44324 6468
rect 43444 3324 43496 3330
rect 43444 3266 43496 3272
rect 44284 480 44312 6462
rect 45468 3324 45520 3330
rect 45468 3266 45520 3272
rect 45480 480 45508 3266
rect 46664 2916 46716 2922
rect 46664 2858 46716 2864
rect 46676 480 46704 2858
rect 47872 480 47900 6886
rect 48964 6588 49016 6594
rect 48964 6530 49016 6536
rect 48976 480 49004 6530
rect 50160 3188 50212 3194
rect 50160 3130 50212 3136
rect 50172 480 50200 3130
rect 50356 2922 50384 279822
rect 51724 275460 51776 275466
rect 51724 275402 51776 275408
rect 51356 5160 51408 5166
rect 51356 5102 51408 5108
rect 50344 2916 50396 2922
rect 50344 2858 50396 2864
rect 51368 480 51396 5102
rect 51736 4010 51764 275402
rect 53116 97986 53144 700470
rect 53194 699816 53250 699825
rect 53194 699751 53250 699760
rect 53208 241466 53236 699751
rect 54484 277024 54536 277030
rect 54484 276966 54536 276972
rect 53196 241460 53248 241466
rect 53196 241402 53248 241408
rect 53104 97980 53156 97986
rect 53104 97922 53156 97928
rect 52552 6656 52604 6662
rect 52552 6598 52604 6604
rect 51724 4004 51776 4010
rect 51724 3946 51776 3952
rect 52564 480 52592 6598
rect 54496 4078 54524 276966
rect 58624 276888 58676 276894
rect 58624 276830 58676 276836
rect 57244 275392 57296 275398
rect 57244 275334 57296 275340
rect 56048 6724 56100 6730
rect 56048 6666 56100 6672
rect 54944 5228 54996 5234
rect 54944 5170 54996 5176
rect 54484 4072 54536 4078
rect 54484 4014 54536 4020
rect 53748 4004 53800 4010
rect 53748 3946 53800 3952
rect 53760 480 53788 3946
rect 54956 480 54984 5170
rect 56060 480 56088 6666
rect 57256 4146 57284 275334
rect 58440 5296 58492 5302
rect 58440 5238 58492 5244
rect 57244 4140 57296 4146
rect 57244 4082 57296 4088
rect 57244 3120 57296 3126
rect 57244 3062 57296 3068
rect 57256 480 57284 3062
rect 58452 480 58480 5238
rect 58636 3398 58664 276830
rect 61384 275324 61436 275330
rect 61384 275266 61436 275272
rect 59636 6792 59688 6798
rect 59636 6734 59688 6740
rect 58624 3392 58676 3398
rect 58624 3334 58676 3340
rect 59648 480 59676 6734
rect 60832 4072 60884 4078
rect 60832 4014 60884 4020
rect 60844 480 60872 4014
rect 61396 3330 61424 275266
rect 65536 189038 65564 701966
rect 68282 699952 68338 699961
rect 68282 699887 68338 699896
rect 68296 255270 68324 699887
rect 68284 255264 68336 255270
rect 68284 255206 68336 255212
rect 65524 189032 65576 189038
rect 65524 188974 65576 188980
rect 71056 150414 71084 702034
rect 72988 700126 73016 703520
rect 79322 701448 79378 701457
rect 79322 701383 79378 701392
rect 72976 700120 73028 700126
rect 72976 700062 73028 700068
rect 79336 346390 79364 701383
rect 89180 700194 89208 703520
rect 105464 700942 105492 703520
rect 105542 701584 105598 701593
rect 105542 701519 105598 701528
rect 105452 700936 105504 700942
rect 105452 700878 105504 700884
rect 89168 700188 89220 700194
rect 89168 700130 89220 700136
rect 79324 346384 79376 346390
rect 79324 346326 79376 346332
rect 105556 293962 105584 701519
rect 137848 701010 137876 703520
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 105544 293956 105596 293962
rect 105544 293898 105596 293904
rect 97264 280152 97316 280158
rect 97264 280094 97316 280100
rect 94504 279200 94556 279206
rect 94504 279142 94556 279148
rect 90364 279132 90416 279138
rect 90364 279074 90416 279080
rect 87604 279064 87656 279070
rect 87604 279006 87656 279012
rect 86224 278996 86276 279002
rect 86224 278938 86276 278944
rect 81348 278248 81400 278254
rect 81348 278190 81400 278196
rect 71044 150408 71096 150414
rect 71044 150350 71096 150356
rect 77392 7880 77444 7886
rect 77392 7822 77444 7828
rect 73804 7812 73856 7818
rect 73804 7754 73856 7760
rect 70308 7676 70360 7682
rect 70308 7618 70360 7624
rect 66720 7608 66772 7614
rect 66720 7550 66772 7556
rect 63224 6860 63276 6866
rect 63224 6802 63276 6808
rect 62028 5364 62080 5370
rect 62028 5306 62080 5312
rect 61384 3324 61436 3330
rect 61384 3266 61436 3272
rect 62040 480 62068 5306
rect 63236 480 63264 6802
rect 65524 5432 65576 5438
rect 65524 5374 65576 5380
rect 64328 2984 64380 2990
rect 64328 2926 64380 2932
rect 64340 480 64368 2926
rect 65536 480 65564 5374
rect 66732 480 66760 7550
rect 69112 5500 69164 5506
rect 69112 5442 69164 5448
rect 67916 4140 67968 4146
rect 67916 4082 67968 4088
rect 67928 480 67956 4082
rect 69124 480 69152 5442
rect 70320 480 70348 7618
rect 72608 4752 72660 4758
rect 72608 4694 72660 4700
rect 71504 3052 71556 3058
rect 71504 2994 71556 3000
rect 71516 480 71544 2994
rect 72620 480 72648 4694
rect 73816 480 73844 7754
rect 76196 4616 76248 4622
rect 76196 4558 76248 4564
rect 75000 3392 75052 3398
rect 75000 3334 75052 3340
rect 75012 480 75040 3334
rect 76208 480 76236 4558
rect 77404 480 77432 7822
rect 79692 4684 79744 4690
rect 79692 4626 79744 4632
rect 78588 2916 78640 2922
rect 78588 2858 78640 2864
rect 78600 480 78628 2858
rect 79704 480 79732 4626
rect 81360 3330 81388 278190
rect 85488 10464 85540 10470
rect 85488 10406 85540 10412
rect 83280 4480 83332 4486
rect 83280 4422 83332 4428
rect 80888 3324 80940 3330
rect 80888 3266 80940 3272
rect 81348 3324 81400 3330
rect 81348 3266 81400 3272
rect 80900 480 80928 3266
rect 82084 3256 82136 3262
rect 82084 3198 82136 3204
rect 82096 480 82124 3198
rect 83292 480 83320 4422
rect 85500 3330 85528 10406
rect 84476 3324 84528 3330
rect 84476 3266 84528 3272
rect 85488 3324 85540 3330
rect 85488 3266 85540 3272
rect 84488 480 84516 3266
rect 86236 3194 86264 278938
rect 86868 4548 86920 4554
rect 86868 4490 86920 4496
rect 86224 3188 86276 3194
rect 86224 3130 86276 3136
rect 85672 3120 85724 3126
rect 85672 3062 85724 3068
rect 85684 480 85712 3062
rect 86880 480 86908 4490
rect 87616 3330 87644 279006
rect 88984 278384 89036 278390
rect 88984 278326 89036 278332
rect 88996 3330 89024 278326
rect 90376 6914 90404 279074
rect 93124 276820 93176 276826
rect 93124 276762 93176 276768
rect 90284 6886 90404 6914
rect 87604 3324 87656 3330
rect 87604 3266 87656 3272
rect 87972 3324 88024 3330
rect 87972 3266 88024 3272
rect 88984 3324 89036 3330
rect 88984 3266 89036 3272
rect 87984 480 88012 3266
rect 89168 2984 89220 2990
rect 89168 2926 89220 2932
rect 89180 480 89208 2926
rect 90284 2922 90312 6886
rect 90364 4412 90416 4418
rect 90364 4354 90416 4360
rect 90272 2916 90324 2922
rect 90272 2858 90324 2864
rect 90376 480 90404 4354
rect 93136 3262 93164 276762
rect 93952 4344 94004 4350
rect 93952 4286 94004 4292
rect 91560 3256 91612 3262
rect 91560 3198 91612 3204
rect 93124 3256 93176 3262
rect 93124 3198 93176 3204
rect 91572 480 91600 3198
rect 93308 3120 93360 3126
rect 93308 3062 93360 3068
rect 93320 2922 93348 3062
rect 92756 2916 92808 2922
rect 92756 2858 92808 2864
rect 93308 2916 93360 2922
rect 93308 2858 93360 2864
rect 92768 480 92796 2858
rect 93964 480 93992 4286
rect 94516 2854 94544 279142
rect 95056 278452 95108 278458
rect 95056 278394 95108 278400
rect 95068 16574 95096 278394
rect 95068 16546 95188 16574
rect 94504 2848 94556 2854
rect 94504 2790 94556 2796
rect 95160 480 95188 16546
rect 97276 2990 97304 280094
rect 111708 280084 111760 280090
rect 111708 280026 111760 280032
rect 101404 280016 101456 280022
rect 101404 279958 101456 279964
rect 99288 278588 99340 278594
rect 99288 278530 99340 278536
rect 97448 4276 97500 4282
rect 97448 4218 97500 4224
rect 97264 2984 97316 2990
rect 97264 2926 97316 2932
rect 96252 2916 96304 2922
rect 96252 2858 96304 2864
rect 96264 480 96292 2858
rect 97460 480 97488 4218
rect 99300 3126 99328 278530
rect 101036 6112 101088 6118
rect 101036 6054 101088 6060
rect 98644 3120 98696 3126
rect 98644 3062 98696 3068
rect 99288 3120 99340 3126
rect 99288 3062 99340 3068
rect 98656 480 98684 3062
rect 99840 2984 99892 2990
rect 99840 2926 99892 2932
rect 99852 480 99880 2926
rect 101048 480 101076 6054
rect 101416 2922 101444 279958
rect 108304 279336 108356 279342
rect 108304 279278 108356 279284
rect 106924 278928 106976 278934
rect 106924 278870 106976 278876
rect 105544 277092 105596 277098
rect 105544 277034 105596 277040
rect 104532 8968 104584 8974
rect 104532 8910 104584 8916
rect 102232 3120 102284 3126
rect 102232 3062 102284 3068
rect 101404 2916 101456 2922
rect 101404 2858 101456 2864
rect 102244 480 102272 3062
rect 103336 2916 103388 2922
rect 103336 2858 103388 2864
rect 103348 480 103376 2858
rect 104544 480 104572 8910
rect 105556 3126 105584 277034
rect 106188 276956 106240 276962
rect 106188 276898 106240 276904
rect 106200 3126 106228 276898
rect 105544 3120 105596 3126
rect 105544 3062 105596 3068
rect 105728 3120 105780 3126
rect 105728 3062 105780 3068
rect 106188 3120 106240 3126
rect 106188 3062 106240 3068
rect 105740 480 105768 3062
rect 106936 3058 106964 278870
rect 108120 9104 108172 9110
rect 108120 9046 108172 9052
rect 106924 3052 106976 3058
rect 106924 2994 106976 3000
rect 106924 2916 106976 2922
rect 106924 2858 106976 2864
rect 106936 480 106964 2858
rect 108132 480 108160 9046
rect 108316 2854 108344 279278
rect 111616 9036 111668 9042
rect 111616 8978 111668 8984
rect 110512 3120 110564 3126
rect 110512 3062 110564 3068
rect 109316 3052 109368 3058
rect 109316 2994 109368 3000
rect 108304 2848 108356 2854
rect 108304 2790 108356 2796
rect 109328 480 109356 2994
rect 110524 480 110552 3062
rect 111628 480 111656 8978
rect 111720 3126 111748 280026
rect 118608 279404 118660 279410
rect 118608 279346 118660 279352
rect 115204 278724 115256 278730
rect 115204 278666 115256 278672
rect 112444 277160 112496 277166
rect 112444 277102 112496 277108
rect 111708 3120 111760 3126
rect 111708 3062 111760 3068
rect 112456 3058 112484 277102
rect 115216 6914 115244 278666
rect 117228 276548 117280 276554
rect 117228 276490 117280 276496
rect 115296 9172 115348 9178
rect 115296 9114 115348 9120
rect 115124 6886 115244 6914
rect 115124 3126 115152 6886
rect 115308 3482 115336 9114
rect 115216 3454 115336 3482
rect 112812 3120 112864 3126
rect 112812 3062 112864 3068
rect 115112 3120 115164 3126
rect 115112 3062 115164 3068
rect 112444 3052 112496 3058
rect 112444 2994 112496 3000
rect 112824 480 112852 3062
rect 114008 3052 114060 3058
rect 114008 2994 114060 3000
rect 114020 480 114048 2994
rect 115216 480 115244 3454
rect 117240 3126 117268 276490
rect 118620 3126 118648 279346
rect 125508 279268 125560 279274
rect 125508 279210 125560 279216
rect 124128 271176 124180 271182
rect 124128 271118 124180 271124
rect 119988 254584 120040 254590
rect 119988 254526 120040 254532
rect 118792 9240 118844 9246
rect 118792 9182 118844 9188
rect 116400 3120 116452 3126
rect 116400 3062 116452 3068
rect 117228 3120 117280 3126
rect 117228 3062 117280 3068
rect 117596 3120 117648 3126
rect 117596 3062 117648 3068
rect 118608 3120 118660 3126
rect 118608 3062 118660 3068
rect 116412 480 116440 3062
rect 117608 480 117636 3062
rect 118804 480 118832 9182
rect 120000 6914 120028 254526
rect 122288 9308 122340 9314
rect 122288 9250 122340 9256
rect 119908 6886 120028 6914
rect 119908 480 119936 6886
rect 121092 2848 121144 2854
rect 121092 2790 121144 2796
rect 121104 480 121132 2790
rect 122300 480 122328 9250
rect 124140 2854 124168 271118
rect 125520 6914 125548 279210
rect 135168 277976 135220 277982
rect 135168 277918 135220 277924
rect 133788 243568 133840 243574
rect 133788 243510 133840 243516
rect 129648 17264 129700 17270
rect 129648 17206 129700 17212
rect 126888 13116 126940 13122
rect 126888 13058 126940 13064
rect 125428 6886 125548 6914
rect 125428 2854 125456 6886
rect 126900 2854 126928 13058
rect 128176 10532 128228 10538
rect 128176 10474 128228 10480
rect 126980 6044 127032 6050
rect 126980 5986 127032 5992
rect 123484 2848 123536 2854
rect 123484 2790 123536 2796
rect 124128 2848 124180 2854
rect 124128 2790 124180 2796
rect 124680 2848 124732 2854
rect 124680 2790 124732 2796
rect 125416 2848 125468 2854
rect 125416 2790 125468 2796
rect 125876 2848 125928 2854
rect 125876 2790 125928 2796
rect 126888 2848 126940 2854
rect 126888 2790 126940 2796
rect 123496 480 123524 2790
rect 124692 480 124720 2790
rect 125888 480 125916 2790
rect 126992 480 127020 5986
rect 128188 480 128216 10474
rect 129660 6914 129688 17206
rect 131764 7948 131816 7954
rect 131764 7890 131816 7896
rect 129384 6886 129688 6914
rect 129384 480 129412 6886
rect 130568 5976 130620 5982
rect 130568 5918 130620 5924
rect 130580 480 130608 5918
rect 131776 480 131804 7890
rect 133800 2854 133828 243510
rect 135180 2854 135208 277918
rect 137928 277364 137980 277370
rect 137928 277306 137980 277312
rect 136456 10736 136508 10742
rect 136456 10678 136508 10684
rect 135260 8016 135312 8022
rect 135260 7958 135312 7964
rect 132960 2848 133012 2854
rect 132960 2790 133012 2796
rect 133788 2848 133840 2854
rect 133788 2790 133840 2796
rect 134156 2848 134208 2854
rect 134156 2790 134208 2796
rect 135168 2848 135220 2854
rect 135168 2790 135220 2796
rect 132972 480 133000 2790
rect 134168 480 134196 2790
rect 135272 480 135300 7958
rect 136468 480 136496 10678
rect 137940 6914 137968 277306
rect 141436 111790 141464 703598
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 330666 703760 330722 703769
rect 330666 703695 330722 703704
rect 148324 702568 148376 702574
rect 148324 702510 148376 702516
rect 144828 277840 144880 277846
rect 144828 277782 144880 277788
rect 141424 111784 141476 111790
rect 141424 111726 141476 111732
rect 142068 71052 142120 71058
rect 142068 70994 142120 71000
rect 140688 10600 140740 10606
rect 140688 10542 140740 10548
rect 138848 9376 138900 9382
rect 138848 9318 138900 9324
rect 137664 6886 137968 6914
rect 137664 480 137692 6886
rect 138860 480 138888 9318
rect 140700 2854 140728 10542
rect 142080 2854 142108 70994
rect 144736 11756 144788 11762
rect 144736 11698 144788 11704
rect 142436 9444 142488 9450
rect 142436 9386 142488 9392
rect 140044 2848 140096 2854
rect 140044 2790 140096 2796
rect 140688 2848 140740 2854
rect 140688 2790 140740 2796
rect 141240 2848 141292 2854
rect 141240 2790 141292 2796
rect 142068 2848 142120 2854
rect 142068 2790 142120 2796
rect 140056 480 140084 2790
rect 141252 480 141280 2790
rect 142448 480 142476 9386
rect 143540 2848 143592 2854
rect 143540 2790 143592 2796
rect 143552 480 143580 2790
rect 144748 480 144776 11698
rect 144840 2854 144868 277782
rect 147588 238060 147640 238066
rect 147588 238002 147640 238008
rect 145932 9512 145984 9518
rect 145932 9454 145984 9460
rect 144828 2848 144880 2854
rect 144828 2790 144880 2796
rect 145944 480 145972 9454
rect 147600 2854 147628 238002
rect 148336 164218 148364 702510
rect 154132 700466 154160 703520
rect 161572 703384 161624 703390
rect 161572 703326 161624 703332
rect 154120 700460 154172 700466
rect 154120 700402 154172 700408
rect 161584 619614 161612 703326
rect 164792 703180 164844 703186
rect 164792 703122 164844 703128
rect 164516 703112 164568 703118
rect 164516 703054 164568 703060
rect 161848 702840 161900 702846
rect 161848 702782 161900 702788
rect 161664 701820 161716 701826
rect 161664 701762 161716 701768
rect 161572 619608 161624 619614
rect 161572 619550 161624 619556
rect 161676 567186 161704 701762
rect 161756 701684 161808 701690
rect 161756 701626 161808 701632
rect 161664 567180 161716 567186
rect 161664 567122 161716 567128
rect 161768 516118 161796 701626
rect 161756 516112 161808 516118
rect 161756 516054 161808 516060
rect 161860 423638 161888 702782
rect 162032 702772 162084 702778
rect 162032 702714 162084 702720
rect 161940 701548 161992 701554
rect 161940 701490 161992 701496
rect 161848 423632 161900 423638
rect 161848 423574 161900 423580
rect 161952 411262 161980 701490
rect 161940 411256 161992 411262
rect 161940 411198 161992 411204
rect 162044 372570 162072 702714
rect 164528 701729 164556 703054
rect 164804 701729 164832 703122
rect 165344 702976 165396 702982
rect 165344 702918 165396 702924
rect 165160 702908 165212 702914
rect 165160 702850 165212 702856
rect 165172 701865 165200 702850
rect 165158 701856 165214 701865
rect 165158 701791 165214 701800
rect 165356 701729 165384 702918
rect 164514 701720 164570 701729
rect 164514 701655 164570 701664
rect 164790 701720 164846 701729
rect 164790 701655 164846 701664
rect 165342 701720 165398 701729
rect 165342 701655 165398 701664
rect 162124 701616 162176 701622
rect 162124 701558 162176 701564
rect 162032 372564 162084 372570
rect 162032 372506 162084 372512
rect 162136 282266 162164 701558
rect 162400 701480 162452 701486
rect 162400 701422 162452 701428
rect 162216 701412 162268 701418
rect 162216 701354 162268 701360
rect 162124 282260 162176 282266
rect 162124 282202 162176 282208
rect 162228 282198 162256 701354
rect 162308 701276 162360 701282
rect 162308 701218 162360 701224
rect 162320 282334 162348 701218
rect 162308 282328 162360 282334
rect 162308 282270 162360 282276
rect 162216 282192 162268 282198
rect 162216 282134 162268 282140
rect 151728 277908 151780 277914
rect 151728 277850 151780 277856
rect 148324 164212 148376 164218
rect 148324 164154 148376 164160
rect 148968 163532 149020 163538
rect 148968 163474 149020 163480
rect 148980 2854 149008 163474
rect 149520 9648 149572 9654
rect 149520 9590 149572 9596
rect 147128 2848 147180 2854
rect 147128 2790 147180 2796
rect 147588 2848 147640 2854
rect 147588 2790 147640 2796
rect 148324 2848 148376 2854
rect 148324 2790 148376 2796
rect 148968 2848 149020 2854
rect 148968 2790 149020 2796
rect 147140 480 147168 2790
rect 148336 480 148364 2790
rect 149532 480 149560 9590
rect 151740 2854 151768 277850
rect 153108 277296 153160 277302
rect 153108 277238 153160 277244
rect 153016 9580 153068 9586
rect 153016 9522 153068 9528
rect 150624 2848 150676 2854
rect 150624 2790 150676 2796
rect 151728 2848 151780 2854
rect 151728 2790 151780 2796
rect 151820 2848 151872 2854
rect 151820 2790 151872 2796
rect 150636 480 150664 2790
rect 151832 480 151860 2790
rect 153028 480 153056 9522
rect 153120 2854 153148 277238
rect 155868 277228 155920 277234
rect 155868 277170 155920 277176
rect 154212 10668 154264 10674
rect 154212 10610 154264 10616
rect 153108 2848 153160 2854
rect 153108 2790 153160 2796
rect 154224 480 154252 10610
rect 155880 2854 155908 277170
rect 160008 276616 160060 276622
rect 160008 276558 160060 276564
rect 158628 11824 158680 11830
rect 158628 11766 158680 11772
rect 156604 8900 156656 8906
rect 156604 8842 156656 8848
rect 155408 2848 155460 2854
rect 155408 2790 155460 2796
rect 155868 2848 155920 2854
rect 155868 2790 155920 2796
rect 155420 480 155448 2790
rect 156616 480 156644 8842
rect 158640 2854 158668 11766
rect 160020 2854 160048 276558
rect 161388 265668 161440 265674
rect 161388 265610 161440 265616
rect 160100 8832 160152 8838
rect 160100 8774 160152 8780
rect 157800 2848 157852 2854
rect 157800 2790 157852 2796
rect 158628 2848 158680 2854
rect 158628 2790 158680 2796
rect 158904 2848 158956 2854
rect 158904 2790 158956 2796
rect 160008 2848 160060 2854
rect 160008 2790 160060 2796
rect 157812 480 157840 2790
rect 158916 480 158944 2790
rect 160112 480 160140 8774
rect 161400 6914 161428 265610
rect 162412 113150 162440 701422
rect 162492 701344 162544 701350
rect 162492 701286 162544 701292
rect 162400 113144 162452 113150
rect 162400 113086 162452 113092
rect 162504 60722 162532 701286
rect 162584 701208 162636 701214
rect 168012 701208 168064 701214
rect 162584 701150 162636 701156
rect 162492 60716 162544 60722
rect 162492 60658 162544 60664
rect 162596 33114 162624 701150
rect 164344 701146 164680 701162
rect 168064 701156 168360 701162
rect 168012 701150 168360 701156
rect 162768 701140 162820 701146
rect 162768 701082 162820 701088
rect 164332 701140 164680 701146
rect 164384 701134 164680 701140
rect 168024 701134 168360 701150
rect 170324 701146 170352 703520
rect 198096 702636 198148 702642
rect 198096 702578 198148 702584
rect 194414 702128 194470 702137
rect 194414 702063 194470 702072
rect 194428 701706 194456 702063
rect 198108 701706 198136 702578
rect 194120 701678 194456 701706
rect 197800 701678 198136 701706
rect 201314 701720 201370 701729
rect 201370 701678 201480 701706
rect 201314 701655 201370 701664
rect 179064 701554 179400 701570
rect 179052 701548 179400 701554
rect 179104 701542 179400 701548
rect 179052 701490 179104 701496
rect 190092 701480 190144 701486
rect 190144 701428 190440 701434
rect 190092 701422 190440 701428
rect 190104 701406 190440 701422
rect 182732 701344 182784 701350
rect 182784 701292 183080 701298
rect 182732 701286 183080 701292
rect 182744 701270 183080 701286
rect 186424 701282 186760 701298
rect 186412 701276 186760 701282
rect 186464 701270 186760 701276
rect 186412 701218 186464 701224
rect 171692 701208 171744 701214
rect 171744 701156 172040 701162
rect 171692 701150 172040 701156
rect 170312 701140 170364 701146
rect 164332 701082 164384 701088
rect 171704 701134 172040 701150
rect 175384 701146 175720 701162
rect 202800 701146 202828 703520
rect 212354 702264 212410 702273
rect 212354 702199 212410 702208
rect 208812 701992 208868 702001
rect 208812 701927 208868 701936
rect 205362 701856 205418 701865
rect 205362 701791 205418 701800
rect 205376 701706 205404 701791
rect 205160 701678 205404 701706
rect 208826 701692 208854 701927
rect 212368 701570 212396 702199
rect 218992 701865 219020 703520
rect 235184 703322 235212 703520
rect 235172 703316 235224 703322
rect 235172 703258 235224 703264
rect 231216 702704 231268 702710
rect 231216 702646 231268 702652
rect 223394 702400 223450 702409
rect 223394 702335 223450 702344
rect 227074 702400 227130 702409
rect 227074 702335 227130 702344
rect 215850 701856 215906 701865
rect 215850 701791 215906 701800
rect 218978 701856 219034 701865
rect 218978 701791 219034 701800
rect 219622 701856 219678 701865
rect 219622 701791 219678 701800
rect 215864 701706 215892 701791
rect 219636 701706 219664 701791
rect 215864 701678 216200 701706
rect 219636 701678 219880 701706
rect 223408 701570 223436 702335
rect 227088 701865 227116 702335
rect 226890 701856 226946 701865
rect 226890 701791 226946 701800
rect 227074 701856 227130 701865
rect 227074 701791 227130 701800
rect 226904 701706 226932 701791
rect 231228 701706 231256 702646
rect 234526 702400 234582 702409
rect 234526 702335 234582 702344
rect 237930 702400 237986 702409
rect 237930 702335 237986 702344
rect 264426 702400 264482 702409
rect 264426 702335 264482 702344
rect 234540 701978 234568 702335
rect 234540 701950 234614 701978
rect 226904 701678 227240 701706
rect 230920 701678 231256 701706
rect 234586 701692 234614 701950
rect 237944 701706 237972 702335
rect 253388 702160 253440 702166
rect 253388 702102 253440 702108
rect 253400 701706 253428 702102
rect 264440 701706 264468 702335
rect 237944 701678 238280 701706
rect 253092 701678 253428 701706
rect 264132 701678 264468 701706
rect 212368 701542 212520 701570
rect 223408 701542 223560 701570
rect 260748 701480 260800 701486
rect 260452 701428 260748 701434
rect 260452 701422 260800 701428
rect 260452 701406 260788 701422
rect 249708 701344 249760 701350
rect 245640 701282 245792 701298
rect 249412 701292 249708 701298
rect 249412 701286 249760 701292
rect 245640 701276 245804 701282
rect 245640 701270 245752 701276
rect 249412 701270 249748 701286
rect 245752 701218 245804 701224
rect 242256 701208 242308 701214
rect 241960 701156 242256 701162
rect 241960 701150 242308 701156
rect 175372 701140 175720 701146
rect 170312 701082 170364 701088
rect 175424 701134 175720 701140
rect 202788 701140 202840 701146
rect 175372 701082 175424 701088
rect 241960 701134 242296 701150
rect 256772 701146 257108 701162
rect 267660 701146 267688 703520
rect 275468 703452 275520 703458
rect 275468 703394 275520 703400
rect 275480 701706 275508 703394
rect 282828 703044 282880 703050
rect 282828 702986 282880 702992
rect 279148 701752 279200 701758
rect 275172 701678 275508 701706
rect 278852 701700 279148 701706
rect 282840 701706 282868 702986
rect 278852 701694 279200 701700
rect 278852 701678 279188 701694
rect 282532 701678 282868 701706
rect 271788 701616 271840 701622
rect 267812 701554 268148 701570
rect 271492 701564 271788 701570
rect 271492 701558 271840 701564
rect 267812 701548 268160 701554
rect 267812 701542 268108 701548
rect 271492 701542 271828 701558
rect 268108 701490 268160 701496
rect 283852 701146 283880 703520
rect 297546 702808 297602 702817
rect 297546 702743 297602 702752
rect 286506 702672 286562 702681
rect 286506 702607 286562 702616
rect 286520 701706 286548 702607
rect 293546 701956 293598 701962
rect 293546 701898 293598 701904
rect 289866 701888 289918 701894
rect 289866 701830 289918 701836
rect 286212 701678 286548 701706
rect 289878 701692 289906 701830
rect 293558 701692 293586 701898
rect 297560 701706 297588 702743
rect 297252 701678 297588 701706
rect 300136 701146 300164 703520
rect 319626 703352 319682 703361
rect 319626 703287 319682 703296
rect 315946 703216 316002 703225
rect 315946 703151 316002 703160
rect 308586 702944 308642 702953
rect 308586 702879 308642 702888
rect 300904 701992 300960 702001
rect 300904 701927 300960 701936
rect 300918 701692 300946 701927
rect 308600 701706 308628 702879
rect 312266 702264 312322 702273
rect 312266 702199 312322 702208
rect 312280 701706 312308 702199
rect 315960 701706 315988 703151
rect 319640 701706 319668 703287
rect 326986 702264 327042 702273
rect 323308 702228 323360 702234
rect 326986 702199 327042 702208
rect 330206 702264 330262 702273
rect 330206 702199 330262 702208
rect 323308 702170 323360 702176
rect 323320 701706 323348 702170
rect 327000 701706 327028 702199
rect 308292 701678 308628 701706
rect 311972 701678 312308 701706
rect 315652 701678 315988 701706
rect 319332 701678 319668 701706
rect 323012 701678 323348 701706
rect 326692 701678 327028 701706
rect 304612 701146 304948 701162
rect 330220 701146 330248 702199
rect 330680 701706 330708 703695
rect 332478 703520 332590 704960
rect 334438 703896 334494 703905
rect 334438 703831 334494 703840
rect 330372 701678 330708 701706
rect 332520 701146 332548 703520
rect 334452 701706 334480 703831
rect 345020 703588 345072 703594
rect 345020 703530 345072 703536
rect 342168 703520 342220 703526
rect 342168 703462 342220 703468
rect 340420 703248 340472 703254
rect 340420 703190 340472 703196
rect 340432 702166 340460 703190
rect 341800 702296 341852 702302
rect 341800 702238 341852 702244
rect 340420 702160 340472 702166
rect 340420 702102 340472 702108
rect 341812 701706 341840 702238
rect 334144 701678 334480 701706
rect 341504 701678 341840 701706
rect 337824 701146 338068 701162
rect 342180 701146 342208 703462
rect 345032 701146 345060 703530
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 396356 703588 396408 703594
rect 396356 703530 396408 703536
rect 346400 703384 346452 703390
rect 346400 703326 346452 703332
rect 346412 702166 346440 703326
rect 348804 702434 348832 703520
rect 362498 703488 362554 703497
rect 351184 703452 351236 703458
rect 351184 703394 351236 703400
rect 352840 703452 352892 703458
rect 362498 703423 362554 703432
rect 352840 703394 352892 703400
rect 349068 703384 349120 703390
rect 349068 703326 349120 703332
rect 348712 702406 348832 702434
rect 346400 702160 346452 702166
rect 346400 702102 346452 702108
rect 345184 701146 345520 701162
rect 348712 701146 348740 702406
rect 349080 701706 349108 703326
rect 350446 702536 350502 702545
rect 350446 702471 350502 702480
rect 350460 702302 350488 702471
rect 351196 702302 351224 703394
rect 350448 702296 350500 702302
rect 350448 702238 350500 702244
rect 351184 702296 351236 702302
rect 351184 702238 351236 702244
rect 352852 701706 352880 703394
rect 358726 702536 358782 702545
rect 356060 702500 356112 702506
rect 358726 702471 358782 702480
rect 361762 702536 361818 702545
rect 361762 702471 361818 702480
rect 356060 702442 356112 702448
rect 348864 701678 349108 701706
rect 352544 701678 352880 701706
rect 356072 701146 356100 702442
rect 358740 702250 358768 702471
rect 358740 702222 359136 702250
rect 358726 702128 358782 702137
rect 358726 702063 358728 702072
rect 358780 702063 358782 702072
rect 358728 702034 358780 702040
rect 359108 702030 359136 702222
rect 360290 702128 360346 702137
rect 360290 702063 360292 702072
rect 360344 702063 360346 702072
rect 360292 702034 360344 702040
rect 361776 702030 361804 702471
rect 362512 702302 362540 703423
rect 364996 702302 365024 703520
rect 385316 703316 385368 703322
rect 385316 703258 385368 703264
rect 367190 702536 367246 702545
rect 367190 702471 367246 702480
rect 374276 702500 374328 702506
rect 367204 702302 367232 702471
rect 374276 702442 374328 702448
rect 362500 702296 362552 702302
rect 362500 702238 362552 702244
rect 363880 702296 363932 702302
rect 363880 702238 363932 702244
rect 364984 702296 365036 702302
rect 364984 702238 365036 702244
rect 367192 702296 367244 702302
rect 367192 702238 367244 702244
rect 359096 702024 359148 702030
rect 359096 701966 359148 701972
rect 361764 702024 361816 702030
rect 361764 701966 361816 701972
rect 363892 701706 363920 702238
rect 363584 701678 363920 701706
rect 374288 701706 374316 702442
rect 385328 701706 385356 703258
rect 392676 702092 392728 702098
rect 392676 702034 392728 702040
rect 392688 701706 392716 702034
rect 396368 701706 396396 703530
rect 397430 703520 397542 704960
rect 407396 703520 407448 703526
rect 413622 703520 413734 704960
rect 418526 703624 418582 703633
rect 418526 703559 418582 703568
rect 374288 701678 374624 701706
rect 385328 701678 385664 701706
rect 392688 701678 393024 701706
rect 396368 701678 396704 701706
rect 356224 701146 356560 701162
rect 359476 701146 359904 701162
rect 367112 701146 367264 701162
rect 370608 701146 370944 701162
rect 378152 701146 378304 701162
rect 381648 701146 381984 701162
rect 389192 701146 389344 701162
rect 397472 701146 397500 703520
rect 407396 703462 407448 703468
rect 407408 701706 407436 703462
rect 407408 701678 407744 701706
rect 400232 701146 400384 701162
rect 403728 701146 404064 701162
rect 411272 701146 411424 701162
rect 413664 701146 413692 703520
rect 418540 701706 418568 703559
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559378 703760 559434 703769
rect 559378 703695 559434 703704
rect 551100 703656 551152 703662
rect 551100 703598 551152 703604
rect 559392 703610 559420 703695
rect 429856 703458 429884 703520
rect 429844 703452 429896 703458
rect 429844 703394 429896 703400
rect 440608 703180 440660 703186
rect 440608 703122 440660 703128
rect 429566 703080 429622 703089
rect 429566 703015 429622 703024
rect 419354 702536 419410 702545
rect 419354 702471 419410 702480
rect 419368 702234 419396 702471
rect 419356 702228 419408 702234
rect 419356 702170 419408 702176
rect 429580 701706 429608 703015
rect 440620 701706 440648 703122
rect 451648 703112 451700 703118
rect 451648 703054 451700 703060
rect 447968 702160 448020 702166
rect 447968 702102 448020 702108
rect 447980 701706 448008 702102
rect 451660 701706 451688 703054
rect 459008 701820 459060 701826
rect 459008 701762 459060 701768
rect 459020 701706 459048 701762
rect 418540 701678 418876 701706
rect 429580 701678 429916 701706
rect 440620 701678 440956 701706
rect 447980 701678 448316 701706
rect 451660 701678 451996 701706
rect 459020 701678 459356 701706
rect 414768 701146 415104 701162
rect 422404 701146 422556 701162
rect 425900 701146 426236 701162
rect 433352 701146 433596 701162
rect 436940 701146 437276 701162
rect 444392 701146 444636 701162
rect 455432 701146 455676 701162
rect 462332 701146 462360 703520
rect 478524 703390 478552 703520
rect 478512 703384 478564 703390
rect 478512 703326 478564 703332
rect 462688 702976 462740 702982
rect 462688 702918 462740 702924
rect 462700 701706 462728 702918
rect 473728 702908 473780 702914
rect 473728 702850 473780 702856
rect 466460 702432 466512 702438
rect 466460 702374 466512 702380
rect 466472 701706 466500 702374
rect 473740 701706 473768 702850
rect 484768 702840 484820 702846
rect 484768 702782 484820 702788
rect 481086 702536 481142 702545
rect 481086 702471 481142 702480
rect 477500 702364 477552 702370
rect 477500 702306 477552 702312
rect 477512 701706 477540 702306
rect 481100 701706 481128 702471
rect 484780 701706 484808 702782
rect 462700 701678 463036 701706
rect 466472 701678 466716 701706
rect 470060 701690 470396 701706
rect 470048 701684 470396 701690
rect 470100 701678 470396 701684
rect 473740 701678 474076 701706
rect 477512 701678 477756 701706
rect 481100 701678 481436 701706
rect 484780 701678 485116 701706
rect 470048 701626 470100 701632
rect 492140 701418 492476 701434
rect 492128 701412 492476 701418
rect 492180 701406 492476 701412
rect 492128 701354 492180 701360
rect 494808 701321 494836 703520
rect 495808 702772 495860 702778
rect 495808 702714 495860 702720
rect 495820 701706 495848 702714
rect 503258 702264 503314 702273
rect 503258 702199 503314 702208
rect 503272 701706 503300 702199
rect 495820 701678 496156 701706
rect 503272 701678 503608 701706
rect 510618 701584 510674 701593
rect 510674 701542 510968 701570
rect 510618 701519 510674 701528
rect 499670 701448 499726 701457
rect 499726 701406 499836 701434
rect 499670 701383 499726 701392
rect 488538 701312 488594 701321
rect 494794 701312 494850 701321
rect 488594 701270 488796 701298
rect 488538 701247 488594 701256
rect 494794 701247 494850 701256
rect 506938 701312 506994 701321
rect 506994 701270 507288 701298
rect 506938 701247 506994 701256
rect 527192 701185 527220 703520
rect 540060 702568 540112 702574
rect 540060 702510 540112 702516
rect 532698 702128 532754 702137
rect 532698 702063 532754 702072
rect 532712 701706 532740 702063
rect 540072 701706 540100 702510
rect 532712 701678 533048 701706
rect 540072 701678 540408 701706
rect 514298 701176 514354 701185
rect 256772 701140 257120 701146
rect 256772 701134 257068 701140
rect 202788 701082 202840 701088
rect 257068 701082 257120 701088
rect 267648 701140 267700 701146
rect 267648 701082 267700 701088
rect 283840 701140 283892 701146
rect 283840 701082 283892 701088
rect 300124 701140 300176 701146
rect 304612 701140 304960 701146
rect 304612 701134 304908 701140
rect 300124 701082 300176 701088
rect 304908 701082 304960 701088
rect 330208 701140 330260 701146
rect 330208 701082 330260 701088
rect 332508 701140 332560 701146
rect 337824 701140 338080 701146
rect 337824 701134 338028 701140
rect 332508 701082 332560 701088
rect 338028 701082 338080 701088
rect 342168 701140 342220 701146
rect 342168 701082 342220 701088
rect 345020 701140 345072 701146
rect 345184 701140 345532 701146
rect 345184 701134 345480 701140
rect 345020 701082 345072 701088
rect 345480 701082 345532 701088
rect 348700 701140 348752 701146
rect 348700 701082 348752 701088
rect 356060 701140 356112 701146
rect 356224 701140 356572 701146
rect 356224 701134 356520 701140
rect 356060 701082 356112 701088
rect 356520 701082 356572 701088
rect 359464 701140 359904 701146
rect 359516 701134 359904 701140
rect 367100 701140 367264 701146
rect 359464 701082 359516 701088
rect 367152 701134 367264 701140
rect 370596 701140 370944 701146
rect 367100 701082 367152 701088
rect 370648 701134 370944 701140
rect 378140 701140 378304 701146
rect 370596 701082 370648 701088
rect 378192 701134 378304 701140
rect 381636 701140 381984 701146
rect 378140 701082 378192 701088
rect 381688 701134 381984 701140
rect 389180 701140 389344 701146
rect 381636 701082 381688 701088
rect 389232 701134 389344 701140
rect 397460 701140 397512 701146
rect 389180 701082 389232 701088
rect 397460 701082 397512 701088
rect 400220 701140 400384 701146
rect 400272 701134 400384 701140
rect 403716 701140 404064 701146
rect 400220 701082 400272 701088
rect 403768 701134 404064 701140
rect 411260 701140 411424 701146
rect 403716 701082 403768 701088
rect 411312 701134 411424 701140
rect 413652 701140 413704 701146
rect 411260 701082 411312 701088
rect 413652 701082 413704 701088
rect 414756 701140 415104 701146
rect 414808 701134 415104 701140
rect 422392 701140 422556 701146
rect 414756 701082 414808 701088
rect 422444 701134 422556 701140
rect 425888 701140 426236 701146
rect 422392 701082 422444 701088
rect 425940 701134 426236 701140
rect 433340 701140 433596 701146
rect 425888 701082 425940 701088
rect 433392 701134 433596 701140
rect 436928 701140 437276 701146
rect 433340 701082 433392 701088
rect 436980 701134 437276 701140
rect 444380 701140 444636 701146
rect 436928 701082 436980 701088
rect 444432 701134 444636 701140
rect 455420 701140 455676 701146
rect 444380 701082 444432 701088
rect 455472 701134 455676 701140
rect 462320 701140 462372 701146
rect 455420 701082 455472 701088
rect 517978 701176 518034 701185
rect 514354 701134 514648 701162
rect 514298 701111 514354 701120
rect 521750 701176 521806 701185
rect 518034 701134 518328 701162
rect 517978 701111 518034 701120
rect 525430 701176 525486 701185
rect 521806 701134 522008 701162
rect 521750 701111 521806 701120
rect 527178 701176 527234 701185
rect 525486 701134 525688 701162
rect 525430 701111 525486 701120
rect 527178 701111 527234 701120
rect 529018 701176 529074 701185
rect 536378 701176 536434 701185
rect 529074 701134 529368 701162
rect 529018 701111 529074 701120
rect 536434 701134 536728 701162
rect 543476 701146 543504 703520
rect 547420 702024 547472 702030
rect 547420 701966 547472 701972
rect 547432 701706 547460 701966
rect 551112 701706 551140 703598
rect 559392 703582 559512 703610
rect 559484 703474 559512 703582
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 559668 703474 559696 703520
rect 559484 703446 559696 703474
rect 577044 703248 577096 703254
rect 577042 703216 577044 703225
rect 577096 703216 577098 703225
rect 577042 703151 577098 703160
rect 576952 703044 577004 703050
rect 576952 702986 577004 702992
rect 576964 702545 576992 702986
rect 576950 702536 577006 702545
rect 576950 702471 577006 702480
rect 583484 701956 583536 701962
rect 583484 701898 583536 701904
rect 582562 701856 582618 701865
rect 562784 701820 562836 701826
rect 582562 701791 582618 701800
rect 562784 701762 562836 701768
rect 562796 701706 562824 701762
rect 547432 701678 547768 701706
rect 551112 701678 551448 701706
rect 555128 701690 555464 701706
rect 555128 701684 555476 701690
rect 555128 701678 555424 701684
rect 562488 701678 562824 701706
rect 582470 701720 582526 701729
rect 582470 701655 582526 701664
rect 555424 701626 555476 701632
rect 566168 701418 566504 701434
rect 566168 701412 566516 701418
rect 566168 701406 566464 701412
rect 566464 701354 566516 701360
rect 573178 701176 573234 701185
rect 543752 701146 544088 701162
rect 558472 701146 558808 701162
rect 543464 701140 543516 701146
rect 536378 701111 536434 701120
rect 462320 701082 462372 701088
rect 543464 701082 543516 701088
rect 543740 701140 544088 701146
rect 543792 701134 544088 701140
rect 558460 701140 558808 701146
rect 543740 701082 543792 701088
rect 558512 701134 558808 701140
rect 569848 701146 570000 701162
rect 569848 701140 570012 701146
rect 569848 701134 569960 701140
rect 558460 701082 558512 701088
rect 580538 701176 580594 701185
rect 573234 701134 573528 701162
rect 577208 701146 577544 701162
rect 577208 701140 577556 701146
rect 577208 701134 577504 701140
rect 573178 701111 573234 701120
rect 569960 701082 570012 701088
rect 580594 701134 580888 701162
rect 580538 701111 580594 701120
rect 577504 701082 577556 701088
rect 162676 701072 162728 701078
rect 162676 701014 162728 701020
rect 162584 33108 162636 33114
rect 162584 33050 162636 33056
rect 162688 20670 162716 701014
rect 162676 20664 162728 20670
rect 162676 20606 162728 20612
rect 162780 10402 162808 701082
rect 582378 700224 582434 700233
rect 582378 700159 582434 700168
rect 580264 282328 580316 282334
rect 580264 282270 580316 282276
rect 162872 281846 163208 281874
rect 163700 281846 164036 281874
rect 164528 281846 164864 281874
rect 162872 278050 162900 281846
rect 163700 278186 163728 281846
rect 164528 278322 164556 281846
rect 165678 281602 165706 281860
rect 165816 281846 166612 281874
rect 167104 281846 167440 281874
rect 167932 281846 168268 281874
rect 168392 281846 169096 281874
rect 169864 281846 170016 281874
rect 170508 281846 170844 281874
rect 171152 281846 171672 281874
rect 172164 281846 172500 281874
rect 173084 281846 173420 281874
rect 173912 281846 174248 281874
rect 174372 281846 175076 281874
rect 175292 281846 175904 281874
rect 176672 281846 176824 281874
rect 176948 281846 177652 281874
rect 178052 281846 178480 281874
rect 178972 281846 179308 281874
rect 179892 281846 180228 281874
rect 180904 281846 181056 281874
rect 181548 281846 181884 281874
rect 182192 281846 182712 281874
rect 165678 281574 165752 281602
rect 164516 278316 164568 278322
rect 164516 278258 164568 278264
rect 163688 278180 163740 278186
rect 163688 278122 163740 278128
rect 162860 278044 162912 278050
rect 162860 277986 162912 277992
rect 165528 10940 165580 10946
rect 165528 10882 165580 10888
rect 162768 10396 162820 10402
rect 162768 10338 162820 10344
rect 163688 8084 163740 8090
rect 163688 8026 163740 8032
rect 161308 6886 161428 6914
rect 161308 480 161336 6886
rect 162492 5908 162544 5914
rect 162492 5850 162544 5856
rect 162504 480 162532 5850
rect 163700 480 163728 8026
rect 165540 3534 165568 10882
rect 165724 6186 165752 281574
rect 165712 6180 165764 6186
rect 165712 6122 165764 6128
rect 164884 3528 164936 3534
rect 164884 3470 164936 3476
rect 165528 3528 165580 3534
rect 165528 3470 165580 3476
rect 164896 480 164924 3470
rect 165816 3466 165844 281846
rect 167104 279478 167132 281846
rect 167092 279472 167144 279478
rect 167092 279414 167144 279420
rect 167932 278526 167960 281846
rect 167920 278520 167972 278526
rect 167920 278462 167972 278468
rect 167184 8220 167236 8226
rect 167184 8162 167236 8168
rect 166080 5840 166132 5846
rect 166080 5782 166132 5788
rect 165804 3460 165856 3466
rect 165804 3402 165856 3408
rect 166092 480 166120 5782
rect 167196 480 167224 8162
rect 168392 6254 168420 281846
rect 169760 279472 169812 279478
rect 169760 279414 169812 279420
rect 169668 11008 169720 11014
rect 169668 10950 169720 10956
rect 168380 6248 168432 6254
rect 168380 6190 168432 6196
rect 169576 6180 169628 6186
rect 169576 6122 169628 6128
rect 168380 3528 168432 3534
rect 168380 3470 168432 3476
rect 168392 480 168420 3470
rect 169588 480 169616 6122
rect 169680 3534 169708 10950
rect 169772 3602 169800 279414
rect 169760 3596 169812 3602
rect 169760 3538 169812 3544
rect 169668 3528 169720 3534
rect 169668 3470 169720 3476
rect 169864 2854 169892 281846
rect 170508 279478 170536 281846
rect 170496 279472 170548 279478
rect 170496 279414 170548 279420
rect 170772 8152 170824 8158
rect 170772 8094 170824 8100
rect 169852 2848 169904 2854
rect 169852 2790 169904 2796
rect 170784 480 170812 8094
rect 171152 4826 171180 281846
rect 172164 278662 172192 281846
rect 173084 279614 173112 281846
rect 173072 279608 173124 279614
rect 173072 279550 173124 279556
rect 173912 279546 173940 281846
rect 173900 279540 173952 279546
rect 173900 279482 173952 279488
rect 172152 278656 172204 278662
rect 172152 278598 172204 278604
rect 174372 277394 174400 281846
rect 174004 277366 174400 277394
rect 171968 8764 172020 8770
rect 171968 8706 172020 8712
rect 171140 4820 171192 4826
rect 171140 4762 171192 4768
rect 171980 480 172008 8706
rect 173164 6248 173216 6254
rect 173164 6190 173216 6196
rect 173176 480 173204 6190
rect 174004 4894 174032 277366
rect 175292 276690 175320 281846
rect 175280 276684 175332 276690
rect 175280 276626 175332 276632
rect 176672 16574 176700 281846
rect 176672 16546 176792 16574
rect 176568 10804 176620 10810
rect 176568 10746 176620 10752
rect 174268 7540 174320 7546
rect 174268 7482 174320 7488
rect 173992 4888 174044 4894
rect 173992 4830 174044 4836
rect 174280 480 174308 7482
rect 176580 3534 176608 10746
rect 176660 5772 176712 5778
rect 176660 5714 176712 5720
rect 175464 3528 175516 3534
rect 175464 3470 175516 3476
rect 176568 3528 176620 3534
rect 176568 3470 176620 3476
rect 175476 480 175504 3470
rect 176672 480 176700 5714
rect 176764 3738 176792 16546
rect 176752 3732 176804 3738
rect 176752 3674 176804 3680
rect 176948 3670 176976 281846
rect 177856 8288 177908 8294
rect 177856 8230 177908 8236
rect 176936 3664 176988 3670
rect 176936 3606 176988 3612
rect 177868 480 177896 8230
rect 178052 4962 178080 281846
rect 178972 277394 179000 281846
rect 179892 279954 179920 281846
rect 179880 279948 179932 279954
rect 179880 279890 179932 279896
rect 180904 279682 180932 281846
rect 180892 279676 180944 279682
rect 180892 279618 180944 279624
rect 180064 279472 180116 279478
rect 180064 279414 180116 279420
rect 178144 277366 179000 277394
rect 178144 276758 178172 277366
rect 178132 276752 178184 276758
rect 178132 276694 178184 276700
rect 179052 10872 179104 10878
rect 179052 10814 179104 10820
rect 178040 4956 178092 4962
rect 178040 4898 178092 4904
rect 179064 480 179092 10814
rect 180076 7750 180104 279414
rect 181548 277394 181576 281846
rect 180904 277366 181576 277394
rect 180064 7744 180116 7750
rect 180064 7686 180116 7692
rect 180248 5704 180300 5710
rect 180248 5646 180300 5652
rect 180260 480 180288 5646
rect 180904 5098 180932 277366
rect 182192 275466 182220 281846
rect 183618 281602 183646 281860
rect 183572 281574 183646 281602
rect 183756 281846 184460 281874
rect 185044 281846 185288 281874
rect 185872 281846 186208 281874
rect 186332 281846 187036 281874
rect 182180 275460 182232 275466
rect 182180 275402 182232 275408
rect 181444 7744 181496 7750
rect 181444 7686 181496 7692
rect 180892 5092 180944 5098
rect 180892 5034 180944 5040
rect 181456 480 181484 7686
rect 183572 3806 183600 281574
rect 183756 6914 183784 281846
rect 185044 277030 185072 281846
rect 185872 279750 185900 281846
rect 185860 279744 185912 279750
rect 185860 279686 185912 279692
rect 185032 277024 185084 277030
rect 185032 276966 185084 276972
rect 184940 7472 184992 7478
rect 184940 7414 184992 7420
rect 183664 6886 183784 6914
rect 183664 5030 183692 6886
rect 183744 5636 183796 5642
rect 183744 5578 183796 5584
rect 183652 5024 183704 5030
rect 183652 4966 183704 4972
rect 183560 3800 183612 3806
rect 183560 3742 183612 3748
rect 182548 3596 182600 3602
rect 182548 3538 182600 3544
rect 182560 480 182588 3538
rect 183756 480 183784 5578
rect 184952 480 184980 7414
rect 186332 6322 186360 281846
rect 187850 281602 187878 281860
rect 187804 281574 187878 281602
rect 188356 281846 188692 281874
rect 189184 281846 189612 281874
rect 190104 281846 190440 281874
rect 190932 281846 191268 281874
rect 191852 281846 192096 281874
rect 192312 281846 193016 281874
rect 193232 281846 193844 281874
rect 187700 279676 187752 279682
rect 187700 279618 187752 279624
rect 186320 6316 186372 6322
rect 186320 6258 186372 6264
rect 187332 6316 187384 6322
rect 187332 6258 187384 6264
rect 186136 3460 186188 3466
rect 186136 3402 186188 3408
rect 186148 480 186176 3402
rect 187344 480 187372 6258
rect 187712 3874 187740 279618
rect 187804 275398 187832 281574
rect 188356 279682 188384 281846
rect 188344 279676 188396 279682
rect 188344 279618 188396 279624
rect 187792 275392 187844 275398
rect 187792 275334 187844 275340
rect 188528 7404 188580 7410
rect 188528 7346 188580 7352
rect 187700 3868 187752 3874
rect 187700 3810 187752 3816
rect 188540 480 188568 7346
rect 189184 6390 189212 281846
rect 190104 279478 190132 281846
rect 190932 279818 190960 281846
rect 190920 279812 190972 279818
rect 190920 279754 190972 279760
rect 191104 279540 191156 279546
rect 191104 279482 191156 279488
rect 190092 279472 190144 279478
rect 190092 279414 190144 279420
rect 189172 6384 189224 6390
rect 189172 6326 189224 6332
rect 190828 6384 190880 6390
rect 190828 6326 190880 6332
rect 189724 3732 189776 3738
rect 189724 3674 189776 3680
rect 189736 480 189764 3674
rect 190840 480 190868 6326
rect 191116 4010 191144 279482
rect 191852 6458 191880 281846
rect 192312 277394 192340 281846
rect 192484 279472 192536 279478
rect 192484 279414 192536 279420
rect 191944 277366 192340 277394
rect 191944 276894 191972 277366
rect 191932 276888 191984 276894
rect 191932 276830 191984 276836
rect 192024 7336 192076 7342
rect 192024 7278 192076 7284
rect 191840 6452 191892 6458
rect 191840 6394 191892 6400
rect 191104 4004 191156 4010
rect 191104 3946 191156 3952
rect 192036 480 192064 7278
rect 192496 4078 192524 279414
rect 192484 4072 192536 4078
rect 192484 4014 192536 4020
rect 193232 3942 193260 281846
rect 194658 281602 194686 281860
rect 194612 281574 194686 281602
rect 194796 281846 195500 281874
rect 196084 281846 196420 281874
rect 196912 281846 197248 281874
rect 197372 281846 198076 281874
rect 198752 281846 198904 281874
rect 199028 281846 199824 281874
rect 200224 281846 200652 281874
rect 201144 281846 201480 281874
rect 201604 281846 202308 281874
rect 202984 281846 203228 281874
rect 203720 281846 204056 281874
rect 204272 281846 204884 281874
rect 194612 6526 194640 281574
rect 194796 275330 194824 281846
rect 196084 279886 196112 281846
rect 196072 279880 196124 279886
rect 196072 279822 196124 279828
rect 196624 279880 196676 279886
rect 196624 279822 196676 279828
rect 195244 279608 195296 279614
rect 195244 279550 195296 279556
rect 194784 275324 194836 275330
rect 194784 275266 194836 275272
rect 194600 6520 194652 6526
rect 194600 6462 194652 6468
rect 194416 6452 194468 6458
rect 194416 6394 194468 6400
rect 193220 3936 193272 3942
rect 193220 3878 193272 3884
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 193232 480 193260 3470
rect 194428 480 194456 6394
rect 195256 4146 195284 279550
rect 195612 7268 195664 7274
rect 195612 7210 195664 7216
rect 195244 4140 195296 4146
rect 195244 4082 195296 4088
rect 195624 480 195652 7210
rect 196636 3398 196664 279822
rect 196912 278118 196940 281846
rect 196900 278112 196952 278118
rect 196900 278054 196952 278060
rect 197372 6594 197400 281846
rect 198752 279002 198780 281846
rect 198740 278996 198792 279002
rect 198740 278938 198792 278944
rect 197360 6588 197412 6594
rect 197360 6530 197412 6536
rect 197912 6520 197964 6526
rect 197912 6462 197964 6468
rect 196808 3800 196860 3806
rect 196808 3742 196860 3748
rect 196624 3392 196676 3398
rect 196624 3334 196676 3340
rect 196820 480 196848 3742
rect 197924 480 197952 6462
rect 199028 5166 199056 281846
rect 199384 279812 199436 279818
rect 199384 279754 199436 279760
rect 199108 7200 199160 7206
rect 199108 7142 199160 7148
rect 199016 5160 199068 5166
rect 199016 5102 199068 5108
rect 199120 480 199148 7142
rect 199396 3330 199424 279754
rect 200224 6662 200252 281846
rect 200764 279676 200816 279682
rect 200764 279618 200816 279624
rect 200212 6656 200264 6662
rect 200212 6598 200264 6604
rect 200304 3664 200356 3670
rect 200304 3606 200356 3612
rect 199384 3324 199436 3330
rect 199384 3266 199436 3272
rect 200316 480 200344 3606
rect 200776 3262 200804 279618
rect 201144 279546 201172 281846
rect 201132 279540 201184 279546
rect 201132 279482 201184 279488
rect 201500 6588 201552 6594
rect 201500 6530 201552 6536
rect 200764 3256 200816 3262
rect 200764 3198 200816 3204
rect 201512 480 201540 6530
rect 201604 5234 201632 281846
rect 202696 7132 202748 7138
rect 202696 7074 202748 7080
rect 201592 5228 201644 5234
rect 201592 5170 201644 5176
rect 202708 480 202736 7074
rect 202984 6730 203012 281846
rect 203524 279540 203576 279546
rect 203524 279482 203576 279488
rect 202972 6724 203024 6730
rect 202972 6666 203024 6672
rect 203536 3194 203564 279482
rect 203720 279070 203748 281846
rect 203708 279064 203760 279070
rect 203708 279006 203760 279012
rect 204272 5302 204300 281846
rect 205698 281602 205726 281860
rect 205652 281574 205726 281602
rect 206296 281846 206632 281874
rect 207032 281846 207460 281874
rect 207584 281846 208288 281874
rect 208872 281846 209208 281874
rect 209792 281846 210036 281874
rect 210252 281846 210864 281874
rect 211356 281846 211692 281874
rect 205652 6798 205680 281574
rect 206296 279478 206324 281846
rect 206284 279472 206336 279478
rect 206284 279414 206336 279420
rect 206376 279472 206428 279478
rect 206376 279414 206428 279420
rect 206388 277394 206416 279414
rect 206296 277366 206416 277394
rect 206192 7064 206244 7070
rect 206192 7006 206244 7012
rect 205640 6792 205692 6798
rect 205640 6734 205692 6740
rect 205088 6656 205140 6662
rect 205088 6598 205140 6604
rect 204260 5296 204312 5302
rect 204260 5238 204312 5244
rect 203892 3868 203944 3874
rect 203892 3810 203944 3816
rect 203524 3188 203576 3194
rect 203524 3130 203576 3136
rect 203904 480 203932 3810
rect 205100 480 205128 6598
rect 206204 480 206232 7006
rect 206296 2990 206324 277366
rect 207032 5370 207060 281846
rect 207584 277394 207612 281846
rect 208492 279744 208544 279750
rect 208492 279686 208544 279692
rect 207124 277366 207612 277394
rect 207124 6866 207152 277366
rect 208504 271182 208532 279686
rect 208872 279138 208900 281846
rect 208860 279132 208912 279138
rect 208860 279074 208912 279080
rect 209044 278520 209096 278526
rect 209044 278462 209096 278468
rect 208492 271176 208544 271182
rect 208492 271118 208544 271124
rect 207112 6860 207164 6866
rect 207112 6802 207164 6808
rect 208584 6724 208636 6730
rect 208584 6666 208636 6672
rect 207020 5364 207072 5370
rect 207020 5306 207072 5312
rect 207388 4072 207440 4078
rect 207388 4014 207440 4020
rect 206284 2984 206336 2990
rect 206284 2926 206336 2932
rect 207400 480 207428 4014
rect 208596 480 208624 6666
rect 209056 3602 209084 278462
rect 209792 5438 209820 281846
rect 210252 277394 210280 281846
rect 211356 279614 211384 281846
rect 212598 281602 212626 281860
rect 212552 281574 212626 281602
rect 212736 281846 213440 281874
rect 213932 281846 214268 281874
rect 214484 281846 215096 281874
rect 215312 281846 216016 281874
rect 216692 281846 216844 281874
rect 216968 281846 217672 281874
rect 218164 281846 218500 281874
rect 219084 281846 219420 281874
rect 219544 281846 220248 281874
rect 220832 281846 221076 281874
rect 221568 281846 221904 281874
rect 222212 281846 222824 281874
rect 211344 279608 211396 279614
rect 211344 279550 211396 279556
rect 209884 277366 210280 277394
rect 209884 7614 209912 277366
rect 209872 7608 209924 7614
rect 209872 7550 209924 7556
rect 212172 6792 212224 6798
rect 212172 6734 212224 6740
rect 209780 5432 209832 5438
rect 209780 5374 209832 5380
rect 209780 5160 209832 5166
rect 209780 5102 209832 5108
rect 209044 3596 209096 3602
rect 209044 3538 209096 3544
rect 209792 480 209820 5102
rect 210976 4004 211028 4010
rect 210976 3946 211028 3952
rect 210988 480 211016 3946
rect 212184 480 212212 6734
rect 212552 5506 212580 281574
rect 212736 7682 212764 281846
rect 213932 278934 213960 281846
rect 213920 278928 213972 278934
rect 213920 278870 213972 278876
rect 214484 277394 214512 281846
rect 214564 279608 214616 279614
rect 214564 279550 214616 279556
rect 214024 277366 214512 277394
rect 212724 7676 212776 7682
rect 212724 7618 212776 7624
rect 212540 5500 212592 5506
rect 212540 5442 212592 5448
rect 214024 4758 214052 277366
rect 214012 4752 214064 4758
rect 214012 4694 214064 4700
rect 214472 4140 214524 4146
rect 214472 4082 214524 4088
rect 213368 3596 213420 3602
rect 213368 3538 213420 3544
rect 213380 480 213408 3538
rect 214484 480 214512 4082
rect 214576 3126 214604 279550
rect 215312 7818 215340 281846
rect 216692 279886 216720 281846
rect 216680 279880 216732 279886
rect 216680 279822 216732 279828
rect 215944 276684 215996 276690
rect 215944 276626 215996 276632
rect 215300 7812 215352 7818
rect 215300 7754 215352 7760
rect 215668 6860 215720 6866
rect 215668 6802 215720 6808
rect 214564 3120 214616 3126
rect 214564 3062 214616 3068
rect 215680 480 215708 6802
rect 215956 3602 215984 276626
rect 216864 5228 216916 5234
rect 216864 5170 216916 5176
rect 215944 3596 215996 3602
rect 215944 3538 215996 3544
rect 216876 480 216904 5170
rect 216968 4622 216996 281846
rect 218164 7886 218192 281846
rect 219084 279206 219112 281846
rect 219072 279200 219124 279206
rect 219072 279142 219124 279148
rect 218152 7880 218204 7886
rect 218152 7822 218204 7828
rect 219544 4690 219572 281846
rect 220832 278254 220860 281846
rect 221464 279880 221516 279886
rect 221464 279822 221516 279828
rect 220820 278248 220872 278254
rect 220820 278190 220872 278196
rect 220728 276888 220780 276894
rect 220728 276830 220780 276836
rect 220740 6914 220768 276830
rect 220464 6886 220768 6914
rect 219532 4684 219584 4690
rect 219532 4626 219584 4632
rect 216956 4616 217008 4622
rect 216956 4558 217008 4564
rect 218060 3936 218112 3942
rect 218060 3878 218112 3884
rect 218072 480 218100 3878
rect 219256 3392 219308 3398
rect 219256 3334 219308 3340
rect 219268 480 219296 3334
rect 220464 480 220492 6886
rect 221476 3058 221504 279822
rect 221568 279818 221596 281846
rect 221740 279880 221792 279886
rect 221740 279822 221792 279828
rect 221556 279812 221608 279818
rect 221556 279754 221608 279760
rect 221752 277394 221780 279822
rect 221568 277366 221780 277394
rect 221568 16574 221596 277366
rect 221568 16546 221688 16574
rect 221556 3596 221608 3602
rect 221556 3538 221608 3544
rect 221464 3052 221516 3058
rect 221464 2994 221516 3000
rect 221568 480 221596 3538
rect 221660 2922 221688 16546
rect 222212 4486 222240 281846
rect 223638 281602 223666 281860
rect 223592 281574 223666 281602
rect 224144 281846 224480 281874
rect 224972 281846 225308 281874
rect 225892 281846 226228 281874
rect 226720 281846 227056 281874
rect 227732 281846 227884 281874
rect 228008 281846 228712 281874
rect 229388 281846 229632 281874
rect 229848 281846 230460 281874
rect 230952 281846 231288 281874
rect 231872 281846 232208 281874
rect 232424 281846 233036 281874
rect 233252 281846 233864 281874
rect 222844 279948 222896 279954
rect 222844 279890 222896 279896
rect 222856 254590 222884 279890
rect 222844 254584 222896 254590
rect 222844 254526 222896 254532
rect 223488 11892 223540 11898
rect 223488 11834 223540 11840
rect 222200 4480 222252 4486
rect 222200 4422 222252 4428
rect 223500 3534 223528 11834
rect 223592 10470 223620 281574
rect 224144 279682 224172 281846
rect 224132 279676 224184 279682
rect 224132 279618 224184 279624
rect 224868 278316 224920 278322
rect 224868 278258 224920 278264
rect 224224 11960 224276 11966
rect 224224 11902 224276 11908
rect 223580 10464 223632 10470
rect 223580 10406 223632 10412
rect 224236 3602 224264 11902
rect 224224 3596 224276 3602
rect 224224 3538 224276 3544
rect 224880 3534 224908 278258
rect 224972 4554 225000 281846
rect 225892 278390 225920 281846
rect 226720 280158 226748 281846
rect 226708 280152 226760 280158
rect 226708 280094 226760 280100
rect 226984 280152 227036 280158
rect 226984 280094 227036 280100
rect 225880 278384 225932 278390
rect 225880 278326 225932 278332
rect 226996 276554 227024 280094
rect 227628 278044 227680 278050
rect 227628 277986 227680 277992
rect 227536 276752 227588 276758
rect 227536 276694 227588 276700
rect 226984 276548 227036 276554
rect 226984 276490 227036 276496
rect 224960 4548 225012 4554
rect 224960 4490 225012 4496
rect 225144 3596 225196 3602
rect 225144 3538 225196 3544
rect 222752 3528 222804 3534
rect 222752 3470 222804 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 223948 3528 224000 3534
rect 223948 3470 224000 3476
rect 224868 3528 224920 3534
rect 224868 3470 224920 3476
rect 221648 2916 221700 2922
rect 221648 2858 221700 2864
rect 222764 480 222792 3470
rect 223960 480 223988 3470
rect 225156 480 225184 3538
rect 226340 3324 226392 3330
rect 226340 3266 226392 3272
rect 226352 480 226380 3266
rect 227548 480 227576 276694
rect 227640 3330 227668 277986
rect 227732 4418 227760 281846
rect 228008 276826 228036 281846
rect 229388 279546 229416 281846
rect 229376 279540 229428 279546
rect 229376 279482 229428 279488
rect 229848 277394 229876 281846
rect 230952 278458 230980 281846
rect 231214 280800 231270 280809
rect 231214 280735 231270 280744
rect 230940 278452 230992 278458
rect 230940 278394 230992 278400
rect 231124 277704 231176 277710
rect 231124 277646 231176 277652
rect 229204 277366 229876 277394
rect 227996 276820 228048 276826
rect 227996 276762 228048 276768
rect 228640 12096 228692 12102
rect 228640 12038 228692 12044
rect 227720 4412 227772 4418
rect 227720 4354 227772 4360
rect 228652 3602 228680 12038
rect 229204 4350 229232 277366
rect 230940 12028 230992 12034
rect 230940 11970 230992 11976
rect 229192 4344 229244 4350
rect 229192 4286 229244 4292
rect 229836 4140 229888 4146
rect 229836 4082 229888 4088
rect 228640 3596 228692 3602
rect 228640 3538 228692 3544
rect 228732 3596 228784 3602
rect 228732 3538 228784 3544
rect 227628 3324 227680 3330
rect 227628 3266 227680 3272
rect 228744 480 228772 3538
rect 229848 480 229876 4082
rect 230952 3602 230980 11970
rect 230940 3596 230992 3602
rect 230940 3538 230992 3544
rect 231032 3596 231084 3602
rect 231032 3538 231084 3544
rect 231044 480 231072 3538
rect 231136 3398 231164 277646
rect 231228 179382 231256 280735
rect 231872 280022 231900 281846
rect 231860 280016 231912 280022
rect 231860 279958 231912 279964
rect 232424 277394 232452 281846
rect 233252 278882 233280 281846
rect 234678 281602 234706 281860
rect 234632 281574 234706 281602
rect 234816 281846 235612 281874
rect 236104 281846 236440 281874
rect 236932 281846 237268 281874
rect 237392 281846 238096 281874
rect 238772 281846 239016 281874
rect 239508 281846 239844 281874
rect 240152 281846 240672 281874
rect 240796 281846 241500 281874
rect 242084 281846 242420 281874
rect 242912 281846 243248 281874
rect 243740 281846 244076 281874
rect 244568 281846 244904 281874
rect 233974 280936 234030 280945
rect 233974 280871 234030 280880
rect 233884 279676 233936 279682
rect 233884 279618 233936 279624
rect 233160 278854 233280 278882
rect 233160 278594 233188 278854
rect 233148 278588 233200 278594
rect 233148 278530 233200 278536
rect 233148 278112 233200 278118
rect 233148 278054 233200 278060
rect 231964 277366 232452 277394
rect 231216 179376 231268 179382
rect 231216 179318 231268 179324
rect 231964 4282 231992 277366
rect 231952 4276 232004 4282
rect 231952 4218 232004 4224
rect 231124 3392 231176 3398
rect 231124 3334 231176 3340
rect 233160 3194 233188 278054
rect 233896 8770 233924 279618
rect 233988 219434 234016 280871
rect 234632 279478 234660 281574
rect 234620 279472 234672 279478
rect 234620 279414 234672 279420
rect 233976 219428 234028 219434
rect 233976 219370 234028 219376
rect 233976 163600 234028 163606
rect 233976 163542 234028 163548
rect 233988 12434 234016 163542
rect 233988 12406 234108 12434
rect 233884 8764 233936 8770
rect 233884 8706 233936 8712
rect 233976 8764 234028 8770
rect 233976 8706 234028 8712
rect 233988 4146 234016 8706
rect 233976 4140 234028 4146
rect 233976 4082 234028 4088
rect 234080 3534 234108 12406
rect 234816 6118 234844 281846
rect 236104 277098 236132 281846
rect 236932 279342 236960 281846
rect 236920 279336 236972 279342
rect 236920 279278 236972 279284
rect 236092 277092 236144 277098
rect 236092 277034 236144 277040
rect 237392 8974 237420 281846
rect 238772 278882 238800 281846
rect 239508 279614 239536 281846
rect 239496 279608 239548 279614
rect 239496 279550 239548 279556
rect 238680 278854 238800 278882
rect 238024 277568 238076 277574
rect 238024 277510 238076 277516
rect 237380 8968 237432 8974
rect 237380 8910 237432 8916
rect 237380 8696 237432 8702
rect 237380 8638 237432 8644
rect 234804 6112 234856 6118
rect 234804 6054 234856 6060
rect 237012 4140 237064 4146
rect 237012 4082 237064 4088
rect 234068 3528 234120 3534
rect 234068 3470 234120 3476
rect 234620 3528 234672 3534
rect 234620 3470 234672 3476
rect 233424 3324 233476 3330
rect 233424 3266 233476 3272
rect 232228 3188 232280 3194
rect 232228 3130 232280 3136
rect 233148 3188 233200 3194
rect 233148 3130 233200 3136
rect 232240 480 232268 3130
rect 233436 480 233464 3266
rect 234632 480 234660 3470
rect 235816 3256 235868 3262
rect 235816 3198 235868 3204
rect 235828 480 235856 3198
rect 237024 480 237052 4082
rect 237392 3398 237420 8638
rect 238036 3466 238064 277510
rect 238680 276962 238708 278854
rect 238668 276956 238720 276962
rect 238668 276898 238720 276904
rect 240152 9110 240180 281846
rect 240796 279698 240824 281846
rect 242084 280090 242112 281846
rect 242072 280084 242124 280090
rect 242072 280026 242124 280032
rect 240244 279670 240824 279698
rect 240244 277166 240272 279670
rect 242808 279608 242860 279614
rect 242808 279550 242860 279556
rect 242716 279472 242768 279478
rect 242716 279414 242768 279420
rect 242164 278248 242216 278254
rect 242164 278190 242216 278196
rect 240784 278180 240836 278186
rect 240784 278122 240836 278128
rect 240232 277160 240284 277166
rect 240232 277102 240284 277108
rect 240140 9104 240192 9110
rect 240140 9046 240192 9052
rect 240140 8968 240192 8974
rect 240140 8910 240192 8916
rect 240152 3534 240180 8910
rect 240796 4078 240824 278122
rect 240784 4072 240836 4078
rect 240784 4014 240836 4020
rect 239312 3528 239364 3534
rect 239312 3470 239364 3476
rect 240140 3528 240192 3534
rect 240140 3470 240192 3476
rect 241704 3528 241756 3534
rect 241704 3470 241756 3476
rect 238024 3460 238076 3466
rect 238024 3402 238076 3408
rect 238116 3460 238168 3466
rect 238116 3402 238168 3408
rect 237380 3392 237432 3398
rect 237380 3334 237432 3340
rect 238128 480 238156 3402
rect 239324 480 239352 3470
rect 240508 3392 240560 3398
rect 240508 3334 240560 3340
rect 240520 480 240548 3334
rect 241716 480 241744 3470
rect 242176 3194 242204 278190
rect 242728 277394 242756 279414
rect 242820 278322 242848 279550
rect 242808 278316 242860 278322
rect 242808 278258 242860 278264
rect 242728 277366 242848 277394
rect 242820 3534 242848 277366
rect 242912 9042 242940 281846
rect 243740 278730 243768 281846
rect 244568 279818 244596 281846
rect 245810 281602 245838 281860
rect 245764 281574 245838 281602
rect 246316 281846 246652 281874
rect 247144 281846 247480 281874
rect 247696 281846 248308 281874
rect 248892 281846 249228 281874
rect 249812 281846 250056 281874
rect 250272 281846 250884 281874
rect 251468 281846 251804 281874
rect 245014 280800 245070 280809
rect 245014 280735 245070 280744
rect 244556 279812 244608 279818
rect 244556 279754 244608 279760
rect 244924 279812 244976 279818
rect 244924 279754 244976 279760
rect 243728 278724 243780 278730
rect 243728 278666 243780 278672
rect 244936 11014 244964 279754
rect 245028 259418 245056 280735
rect 245016 259412 245068 259418
rect 245016 259354 245068 259360
rect 245016 12164 245068 12170
rect 245016 12106 245068 12112
rect 244924 11008 244976 11014
rect 244924 10950 244976 10956
rect 242900 9036 242952 9042
rect 242900 8978 242952 8984
rect 242900 4820 242952 4826
rect 242900 4762 242952 4768
rect 242808 3528 242860 3534
rect 242808 3470 242860 3476
rect 242164 3188 242216 3194
rect 242164 3130 242216 3136
rect 242912 480 242940 4762
rect 245028 3262 245056 12106
rect 245764 9178 245792 281574
rect 246316 280158 246344 281846
rect 246304 280152 246356 280158
rect 246304 280094 246356 280100
rect 247144 279410 247172 281846
rect 247132 279404 247184 279410
rect 247132 279346 247184 279352
rect 246304 277772 246356 277778
rect 246304 277714 246356 277720
rect 245752 9172 245804 9178
rect 245752 9114 245804 9120
rect 246316 3670 246344 277714
rect 247696 277394 247724 281846
rect 248892 279954 248920 281846
rect 248880 279948 248932 279954
rect 248880 279890 248932 279896
rect 249064 279948 249116 279954
rect 249064 279890 249116 279896
rect 247144 277366 247724 277394
rect 247144 9246 247172 277366
rect 249076 10742 249104 279890
rect 249812 279886 249840 281846
rect 249800 279880 249852 279886
rect 249800 279822 249852 279828
rect 249708 279404 249760 279410
rect 249708 279346 249760 279352
rect 249064 10736 249116 10742
rect 249064 10678 249116 10684
rect 247132 9240 247184 9246
rect 247132 9182 247184 9188
rect 246396 4888 246448 4894
rect 246396 4830 246448 4836
rect 246304 3664 246356 3670
rect 246304 3606 246356 3612
rect 245200 3528 245252 3534
rect 245200 3470 245252 3476
rect 245016 3256 245068 3262
rect 245016 3198 245068 3204
rect 244096 3120 244148 3126
rect 244096 3062 244148 3068
rect 244108 480 244136 3062
rect 245212 480 245240 3470
rect 246408 480 246436 4830
rect 247592 4072 247644 4078
rect 247592 4014 247644 4020
rect 247604 480 247632 4014
rect 249720 3670 249748 279346
rect 250272 277394 250300 281846
rect 251468 279750 251496 281846
rect 252618 281602 252646 281860
rect 252572 281574 252646 281602
rect 252756 281846 253460 281874
rect 254044 281846 254288 281874
rect 254872 281846 255208 281874
rect 255332 281846 256036 281874
rect 256712 281846 256864 281874
rect 256988 281846 257692 281874
rect 258092 281846 258612 281874
rect 259104 281846 259440 281874
rect 259564 281846 260268 281874
rect 260852 281846 261096 281874
rect 261680 281846 262016 281874
rect 262232 281846 262844 281874
rect 252008 279880 252060 279886
rect 252008 279822 252060 279828
rect 251456 279744 251508 279750
rect 251456 279686 251508 279692
rect 251824 279744 251876 279750
rect 251824 279686 251876 279692
rect 250444 277636 250496 277642
rect 250444 277578 250496 277584
rect 249904 277366 250300 277394
rect 249904 9314 249932 277366
rect 249892 9308 249944 9314
rect 249892 9250 249944 9256
rect 250456 4010 250484 277578
rect 251836 10538 251864 279686
rect 251916 279540 251968 279546
rect 251916 279482 251968 279488
rect 251928 10946 251956 279482
rect 252020 265674 252048 279822
rect 252572 279274 252600 281574
rect 252560 279268 252612 279274
rect 252560 279210 252612 279216
rect 252008 265668 252060 265674
rect 252008 265610 252060 265616
rect 252756 13122 252784 281846
rect 253204 277432 253256 277438
rect 253204 277374 253256 277380
rect 252744 13116 252796 13122
rect 252744 13058 252796 13064
rect 251916 10940 251968 10946
rect 251916 10882 251968 10888
rect 251824 10532 251876 10538
rect 251824 10474 251876 10480
rect 252008 10532 252060 10538
rect 252008 10474 252060 10480
rect 250444 4004 250496 4010
rect 250444 3946 250496 3952
rect 252020 3874 252048 10474
rect 252008 3868 252060 3874
rect 252008 3810 252060 3816
rect 253216 3738 253244 277374
rect 254044 6050 254072 281846
rect 254872 279750 254900 281846
rect 254860 279744 254912 279750
rect 254860 279686 254912 279692
rect 255332 17270 255360 281846
rect 255412 280084 255464 280090
rect 255412 280026 255464 280032
rect 255424 277370 255452 280026
rect 255412 277364 255464 277370
rect 255412 277306 255464 277312
rect 255964 36576 256016 36582
rect 255964 36518 256016 36524
rect 255320 17264 255372 17270
rect 255320 17206 255372 17212
rect 254032 6044 254084 6050
rect 254032 5986 254084 5992
rect 253480 4956 253532 4962
rect 253480 4898 253532 4904
rect 253204 3732 253256 3738
rect 253204 3674 253256 3680
rect 248788 3664 248840 3670
rect 248788 3606 248840 3612
rect 249708 3664 249760 3670
rect 249708 3606 249760 3612
rect 252376 3664 252428 3670
rect 252376 3606 252428 3612
rect 248800 480 248828 3606
rect 249984 3188 250036 3194
rect 249984 3130 250036 3136
rect 249996 480 250024 3130
rect 251180 3052 251232 3058
rect 251180 2994 251232 3000
rect 251192 480 251220 2994
rect 252388 480 252416 3606
rect 253492 480 253520 4898
rect 254676 3868 254728 3874
rect 254676 3810 254728 3816
rect 254688 480 254716 3810
rect 255976 3806 256004 36518
rect 256712 5982 256740 281846
rect 256988 7954 257016 281846
rect 258092 243574 258120 281846
rect 258724 278384 258776 278390
rect 258724 278326 258776 278332
rect 258080 243568 258132 243574
rect 258080 243510 258132 243516
rect 258080 9104 258132 9110
rect 258080 9046 258132 9052
rect 256976 7948 257028 7954
rect 256976 7890 257028 7896
rect 256700 5976 256752 5982
rect 256700 5918 256752 5924
rect 257068 5092 257120 5098
rect 257068 5034 257120 5040
rect 255964 3800 256016 3806
rect 255964 3742 256016 3748
rect 255872 3256 255924 3262
rect 255872 3198 255924 3204
rect 255884 480 255912 3198
rect 257080 480 257108 5034
rect 258092 3194 258120 9046
rect 258172 4004 258224 4010
rect 258172 3946 258224 3952
rect 258184 3330 258212 3946
rect 258172 3324 258224 3330
rect 258172 3266 258224 3272
rect 258264 3324 258316 3330
rect 258264 3266 258316 3272
rect 258080 3188 258132 3194
rect 258080 3130 258132 3136
rect 258276 480 258304 3266
rect 258736 3058 258764 278326
rect 259104 277982 259132 281846
rect 259092 277976 259144 277982
rect 259092 277918 259144 277924
rect 258816 243568 258868 243574
rect 258816 243510 258868 243516
rect 258828 4010 258856 243510
rect 259564 8022 259592 281846
rect 260852 279954 260880 281846
rect 261680 280090 261708 281846
rect 261668 280084 261720 280090
rect 261668 280026 261720 280032
rect 260840 279948 260892 279954
rect 260840 279890 260892 279896
rect 260104 278316 260156 278322
rect 260104 278258 260156 278264
rect 259552 8016 259604 8022
rect 259552 7958 259604 7964
rect 258816 4004 258868 4010
rect 258816 3946 258868 3952
rect 259460 3732 259512 3738
rect 259460 3674 259512 3680
rect 258724 3052 258776 3058
rect 258724 2994 258776 3000
rect 259472 480 259500 3674
rect 260116 3330 260144 278258
rect 262232 9382 262260 281846
rect 263658 281602 263686 281860
rect 263612 281574 263686 281602
rect 263796 281846 264500 281874
rect 265084 281846 265420 281874
rect 265912 281846 266248 281874
rect 266372 281846 267076 281874
rect 267752 281846 267904 281874
rect 268028 281846 268824 281874
rect 269224 281846 269652 281874
rect 270144 281846 270480 281874
rect 270972 281846 271308 281874
rect 271892 281846 272228 281874
rect 272720 281846 273056 281874
rect 273272 281846 273884 281874
rect 274652 281846 274804 281874
rect 274928 281846 275632 281874
rect 276032 281846 276460 281874
rect 276584 281846 277288 281874
rect 277412 281846 278208 281874
rect 278792 281846 279036 281874
rect 279252 281846 279864 281874
rect 280172 281846 280692 281874
rect 262312 278860 262364 278866
rect 262312 278802 262364 278808
rect 262324 277846 262352 278802
rect 262312 277840 262364 277846
rect 262312 277782 262364 277788
rect 262864 277500 262916 277506
rect 262864 277442 262916 277448
rect 262220 9376 262272 9382
rect 262220 9318 262272 9324
rect 260656 5024 260708 5030
rect 260656 4966 260708 4972
rect 260104 3324 260156 3330
rect 260104 3266 260156 3272
rect 260668 480 260696 4966
rect 262876 3942 262904 277442
rect 263612 10606 263640 281574
rect 263796 71058 263824 281846
rect 263784 71052 263836 71058
rect 263784 70994 263836 71000
rect 263600 10600 263652 10606
rect 263600 10542 263652 10548
rect 265084 9450 265112 281846
rect 265912 278866 265940 281846
rect 265900 278860 265952 278866
rect 265900 278802 265952 278808
rect 266372 11762 266400 281846
rect 267004 277160 267056 277166
rect 267004 277102 267056 277108
rect 266360 11756 266412 11762
rect 266360 11698 266412 11704
rect 265072 9444 265124 9450
rect 265072 9386 265124 9392
rect 264152 9036 264204 9042
rect 264152 8978 264204 8984
rect 262864 3936 262916 3942
rect 262864 3878 262916 3884
rect 261760 3868 261812 3874
rect 261760 3810 261812 3816
rect 261772 480 261800 3810
rect 262956 3188 263008 3194
rect 262956 3130 263008 3136
rect 262968 480 262996 3130
rect 264164 480 264192 8978
rect 265348 4004 265400 4010
rect 265348 3946 265400 3952
rect 265360 480 265388 3946
rect 266544 3936 266596 3942
rect 266544 3878 266596 3884
rect 266556 480 266584 3878
rect 267016 3126 267044 277102
rect 267752 9518 267780 281846
rect 268028 238066 268056 281846
rect 269120 279404 269172 279410
rect 269120 279346 269172 279352
rect 268016 238060 268068 238066
rect 268016 238002 268068 238008
rect 268384 10464 268436 10470
rect 268384 10406 268436 10412
rect 267740 9512 267792 9518
rect 267740 9454 267792 9460
rect 267832 9240 267884 9246
rect 267832 9182 267884 9188
rect 267844 3398 267872 9182
rect 268396 4010 268424 10406
rect 269132 9654 269160 279346
rect 269224 163538 269252 281846
rect 270144 279410 270172 281846
rect 270132 279404 270184 279410
rect 270132 279346 270184 279352
rect 270972 277914 271000 281846
rect 271892 279698 271920 281846
rect 271800 279670 271920 279698
rect 271144 278452 271196 278458
rect 271144 278394 271196 278400
rect 270960 277908 271012 277914
rect 270960 277850 271012 277856
rect 269212 163532 269264 163538
rect 269212 163474 269264 163480
rect 269120 9648 269172 9654
rect 269120 9590 269172 9596
rect 269120 9172 269172 9178
rect 269120 9114 269172 9120
rect 268384 4004 268436 4010
rect 268384 3946 268436 3952
rect 269132 3806 269160 9114
rect 269120 3800 269172 3806
rect 269120 3742 269172 3748
rect 267832 3392 267884 3398
rect 267832 3334 267884 3340
rect 270040 3392 270092 3398
rect 270040 3334 270092 3340
rect 267004 3120 267056 3126
rect 267004 3062 267056 3068
rect 268844 3120 268896 3126
rect 268844 3062 268896 3068
rect 267740 2984 267792 2990
rect 267740 2926 267792 2932
rect 267752 480 267780 2926
rect 268856 480 268884 3062
rect 270052 480 270080 3334
rect 271156 2990 271184 278394
rect 271800 277302 271828 279670
rect 272720 277394 272748 281846
rect 271984 277366 272748 277394
rect 271788 277296 271840 277302
rect 271788 277238 271840 277244
rect 271984 9586 272012 277366
rect 273272 10674 273300 281846
rect 274652 279698 274680 281846
rect 274560 279670 274680 279698
rect 273904 277296 273956 277302
rect 273904 277238 273956 277244
rect 273260 10668 273312 10674
rect 273260 10610 273312 10616
rect 271972 9580 272024 9586
rect 271972 9522 272024 9528
rect 271236 6112 271288 6118
rect 271236 6054 271288 6060
rect 271144 2984 271196 2990
rect 271144 2926 271196 2932
rect 271248 480 271276 6054
rect 273916 4078 273944 277238
rect 274560 277234 274588 279670
rect 274548 277228 274600 277234
rect 274548 277170 274600 277176
rect 274928 8906 274956 281846
rect 276032 11830 276060 281846
rect 276584 277394 276612 281846
rect 276664 279948 276716 279954
rect 276664 279890 276716 279896
rect 276124 277366 276612 277394
rect 276124 276622 276152 277366
rect 276112 276616 276164 276622
rect 276112 276558 276164 276564
rect 276020 11824 276072 11830
rect 276020 11766 276072 11772
rect 274916 8900 274968 8906
rect 274916 8842 274968 8848
rect 274824 6044 274876 6050
rect 274824 5986 274876 5992
rect 273904 4072 273956 4078
rect 273904 4014 273956 4020
rect 272432 4004 272484 4010
rect 272432 3946 272484 3952
rect 272444 480 272472 3946
rect 273628 3800 273680 3806
rect 273628 3742 273680 3748
rect 273640 480 273668 3742
rect 274836 480 274864 5986
rect 276676 5234 276704 279890
rect 277412 8838 277440 281846
rect 278792 279886 278820 281846
rect 278780 279880 278832 279886
rect 278780 279822 278832 279828
rect 278044 278724 278096 278730
rect 278044 278666 278096 278672
rect 277400 8832 277452 8838
rect 277400 8774 277452 8780
rect 276664 5228 276716 5234
rect 276664 5170 276716 5176
rect 278056 3874 278084 278666
rect 279252 277394 279280 281846
rect 278884 277366 279280 277394
rect 278320 5976 278372 5982
rect 278320 5918 278372 5924
rect 278044 3868 278096 3874
rect 278044 3810 278096 3816
rect 277124 3324 277176 3330
rect 277124 3266 277176 3272
rect 276020 3052 276072 3058
rect 276020 2994 276072 3000
rect 276032 480 276060 2994
rect 277136 480 277164 3266
rect 278332 480 278360 5918
rect 278884 5914 278912 277366
rect 280172 8090 280200 281846
rect 281598 281602 281626 281860
rect 281552 281574 281626 281602
rect 281736 281846 282440 281874
rect 283024 281846 283268 281874
rect 283760 281846 284096 281874
rect 284312 281846 285016 281874
rect 281552 279750 281580 281574
rect 281540 279744 281592 279750
rect 281540 279686 281592 279692
rect 280804 277092 280856 277098
rect 280804 277034 280856 277040
rect 280160 8084 280212 8090
rect 280160 8026 280212 8032
rect 278872 5908 278924 5914
rect 278872 5850 278924 5856
rect 280712 4072 280764 4078
rect 280712 4014 280764 4020
rect 279516 3868 279568 3874
rect 279516 3810 279568 3816
rect 279528 480 279556 3810
rect 280724 480 280752 4014
rect 280816 3126 280844 277034
rect 281736 5846 281764 281846
rect 282184 276820 282236 276826
rect 282184 276762 282236 276768
rect 281724 5840 281776 5846
rect 281724 5782 281776 5788
rect 281908 5228 281960 5234
rect 281908 5170 281960 5176
rect 280804 3120 280856 3126
rect 280804 3062 280856 3068
rect 281920 480 281948 5170
rect 282196 4010 282224 276762
rect 283024 8226 283052 281846
rect 283760 279818 283788 281846
rect 283748 279812 283800 279818
rect 283748 279754 283800 279760
rect 283012 8220 283064 8226
rect 283012 8162 283064 8168
rect 284312 6186 284340 281846
rect 285830 281602 285858 281860
rect 285784 281574 285858 281602
rect 286336 281846 286672 281874
rect 287072 281846 287500 281874
rect 287624 281846 288420 281874
rect 288544 281846 289248 281874
rect 289832 281846 290076 281874
rect 290568 281846 290904 281874
rect 291212 281846 291824 281874
rect 284944 277024 284996 277030
rect 284944 276966 284996 276972
rect 284300 6180 284352 6186
rect 284300 6122 284352 6128
rect 282184 4004 282236 4010
rect 282184 3946 282236 3952
rect 283104 4004 283156 4010
rect 283104 3946 283156 3952
rect 283116 480 283144 3946
rect 284300 3120 284352 3126
rect 284300 3062 284352 3068
rect 284312 480 284340 3062
rect 284956 3058 284984 276966
rect 285784 8158 285812 281574
rect 286336 279682 286364 281846
rect 286324 279676 286376 279682
rect 286324 279618 286376 279624
rect 286324 276956 286376 276962
rect 286324 276898 286376 276904
rect 285772 8152 285824 8158
rect 285772 8094 285824 8100
rect 285404 5296 285456 5302
rect 285404 5238 285456 5244
rect 284944 3052 284996 3058
rect 284944 2994 284996 3000
rect 285416 480 285444 5238
rect 286336 3874 286364 276898
rect 287072 6254 287100 281846
rect 287624 277394 287652 281846
rect 287164 277366 287652 277394
rect 287164 7546 287192 277366
rect 288544 10810 288572 281846
rect 289084 278588 289136 278594
rect 289084 278530 289136 278536
rect 288532 10804 288584 10810
rect 288532 10746 288584 10752
rect 287152 7540 287204 7546
rect 287152 7482 287204 7488
rect 287060 6248 287112 6254
rect 287060 6190 287112 6196
rect 288992 5364 289044 5370
rect 288992 5306 289044 5312
rect 287796 4072 287848 4078
rect 287796 4014 287848 4020
rect 286324 3868 286376 3874
rect 286324 3810 286376 3816
rect 286600 3052 286652 3058
rect 286600 2994 286652 3000
rect 286612 480 286640 2994
rect 287808 480 287836 4014
rect 289004 480 289032 5306
rect 289096 3058 289124 278530
rect 289832 5778 289860 281846
rect 290568 277394 290596 281846
rect 289924 277366 290596 277394
rect 289924 8294 289952 277366
rect 291212 10878 291240 281846
rect 292638 281602 292666 281860
rect 292592 281574 292666 281602
rect 292776 281846 293480 281874
rect 293972 281846 294308 281874
rect 294524 281846 295228 281874
rect 295352 281846 296056 281874
rect 296732 281846 296884 281874
rect 297008 281846 297804 281874
rect 298112 281846 298632 281874
rect 299124 281846 299460 281874
rect 299584 281846 300288 281874
rect 300872 281846 301208 281874
rect 301700 281846 302036 281874
rect 302252 281846 302864 281874
rect 291844 278656 291896 278662
rect 291844 278598 291896 278604
rect 291200 10872 291252 10878
rect 291200 10814 291252 10820
rect 289912 8288 289964 8294
rect 289912 8230 289964 8236
rect 291856 6914 291884 278598
rect 292488 7608 292540 7614
rect 292488 7550 292540 7556
rect 291304 6886 291884 6914
rect 289820 5772 289872 5778
rect 289820 5714 289872 5720
rect 291304 4010 291332 6886
rect 291292 4004 291344 4010
rect 291292 3946 291344 3952
rect 291384 4004 291436 4010
rect 291384 3946 291436 3952
rect 289084 3052 289136 3058
rect 289084 2994 289136 3000
rect 290188 3052 290240 3058
rect 290188 2994 290240 3000
rect 290200 480 290228 2994
rect 291396 480 291424 3946
rect 292500 3058 292528 7550
rect 292592 5710 292620 281574
rect 292776 7750 292804 281846
rect 293224 279676 293276 279682
rect 293224 279618 293276 279624
rect 292764 7744 292816 7750
rect 292764 7686 292816 7692
rect 292580 5704 292632 5710
rect 292580 5646 292632 5652
rect 292580 5432 292632 5438
rect 292580 5374 292632 5380
rect 292488 3052 292540 3058
rect 292488 2994 292540 3000
rect 292592 480 292620 5374
rect 293236 4010 293264 279618
rect 293972 278526 294000 281846
rect 293960 278520 294012 278526
rect 293960 278462 294012 278468
rect 294524 277394 294552 281846
rect 293972 277366 294552 277394
rect 293972 5642 294000 277366
rect 295352 7478 295380 281846
rect 295984 280016 296036 280022
rect 295984 279958 296036 279964
rect 295340 7472 295392 7478
rect 295340 7414 295392 7420
rect 293960 5636 294012 5642
rect 293960 5578 294012 5584
rect 295996 5166 296024 279958
rect 296732 277710 296760 281846
rect 296720 277704 296772 277710
rect 296720 277646 296772 277652
rect 297008 277394 297036 281846
rect 296732 277366 297036 277394
rect 296732 6322 296760 277366
rect 298112 7410 298140 281846
rect 299124 277438 299152 281846
rect 299388 279744 299440 279750
rect 299388 279686 299440 279692
rect 299112 277432 299164 277438
rect 299112 277374 299164 277380
rect 298376 7676 298428 7682
rect 298376 7618 298428 7624
rect 298100 7404 298152 7410
rect 298100 7346 298152 7352
rect 296720 6316 296772 6322
rect 296720 6258 296772 6264
rect 295984 5160 296036 5166
rect 295984 5102 296036 5108
rect 296076 5160 296128 5166
rect 296076 5102 296128 5108
rect 294880 4072 294932 4078
rect 294880 4014 294932 4020
rect 293224 4004 293276 4010
rect 293224 3946 293276 3952
rect 293684 3052 293736 3058
rect 293684 2994 293736 3000
rect 293696 480 293724 2994
rect 294892 480 294920 4014
rect 296088 480 296116 5102
rect 298388 2990 298416 7618
rect 299400 3398 299428 279686
rect 299584 6390 299612 281846
rect 300124 279404 300176 279410
rect 300124 279346 300176 279352
rect 299572 6384 299624 6390
rect 299572 6326 299624 6332
rect 299664 4752 299716 4758
rect 299664 4694 299716 4700
rect 298468 3392 298520 3398
rect 298468 3334 298520 3340
rect 299388 3392 299440 3398
rect 299388 3334 299440 3340
rect 297272 2984 297324 2990
rect 297272 2926 297324 2932
rect 298376 2984 298428 2990
rect 298376 2926 298428 2932
rect 297284 480 297312 2926
rect 298480 480 298508 3334
rect 299676 480 299704 4694
rect 300136 3126 300164 279346
rect 300872 7342 300900 281846
rect 301700 277574 301728 281846
rect 301688 277568 301740 277574
rect 301688 277510 301740 277516
rect 300860 7336 300912 7342
rect 300860 7278 300912 7284
rect 302252 6458 302280 281846
rect 303678 281602 303706 281860
rect 303632 281574 303706 281602
rect 303816 281846 304612 281874
rect 305012 281846 305440 281874
rect 305748 281846 306268 281874
rect 306392 281846 307096 281874
rect 307772 281846 308016 281874
rect 308232 281846 308844 281874
rect 309244 281846 309672 281874
rect 310164 281846 310500 281874
rect 310624 281846 311420 281874
rect 311912 281846 312248 281874
rect 312372 281846 313076 281874
rect 313568 281846 313904 281874
rect 314672 281846 314824 281874
rect 314948 281846 315652 281874
rect 316144 281846 316480 281874
rect 316972 281846 317308 281874
rect 317432 281846 318228 281874
rect 318812 281846 319056 281874
rect 319548 281846 319884 281874
rect 320192 281846 320804 281874
rect 302884 280084 302936 280090
rect 302884 280026 302936 280032
rect 302240 6452 302292 6458
rect 302240 6394 302292 6400
rect 300124 3120 300176 3126
rect 300124 3062 300176 3068
rect 300768 2984 300820 2990
rect 300768 2926 300820 2932
rect 300780 480 300808 2926
rect 301964 2916 302016 2922
rect 301964 2858 302016 2864
rect 301976 480 302004 2858
rect 302896 2854 302924 280026
rect 303632 7274 303660 281574
rect 303816 36582 303844 281846
rect 303804 36576 303856 36582
rect 303804 36518 303856 36524
rect 304356 7744 304408 7750
rect 304356 7686 304408 7692
rect 303620 7268 303672 7274
rect 303620 7210 303672 7216
rect 303160 5500 303212 5506
rect 303160 5442 303212 5448
rect 302884 2848 302936 2854
rect 302884 2790 302936 2796
rect 303172 480 303200 5442
rect 304368 480 304396 7686
rect 305012 6526 305040 281846
rect 305748 277394 305776 281846
rect 306288 279812 306340 279818
rect 306288 279754 306340 279760
rect 305104 277366 305776 277394
rect 305104 7206 305132 277366
rect 305092 7200 305144 7206
rect 305092 7142 305144 7148
rect 305000 6520 305052 6526
rect 305000 6462 305052 6468
rect 306300 3398 306328 279754
rect 306392 12170 306420 281846
rect 307024 279268 307076 279274
rect 307024 279210 307076 279216
rect 306380 12164 306432 12170
rect 306380 12106 306432 12112
rect 306748 4684 306800 4690
rect 306748 4626 306800 4632
rect 305552 3392 305604 3398
rect 305552 3334 305604 3340
rect 306288 3392 306340 3398
rect 306288 3334 306340 3340
rect 305564 480 305592 3334
rect 306760 480 306788 4626
rect 307036 3330 307064 279210
rect 307772 6594 307800 281846
rect 308232 277394 308260 281846
rect 309140 279880 309192 279886
rect 309140 279822 309192 279828
rect 307864 277366 308260 277394
rect 307864 7138 307892 277366
rect 307852 7132 307904 7138
rect 307852 7074 307904 7080
rect 309152 6662 309180 279822
rect 309244 10538 309272 281846
rect 310164 279886 310192 281846
rect 310152 279880 310204 279886
rect 310152 279822 310204 279828
rect 309232 10532 309284 10538
rect 309232 10474 309284 10480
rect 310624 7070 310652 281846
rect 311912 277778 311940 281846
rect 311900 277772 311952 277778
rect 311900 277714 311952 277720
rect 312372 277394 312400 281846
rect 313568 280022 313596 281846
rect 313556 280016 313608 280022
rect 313556 279958 313608 279964
rect 313188 279880 313240 279886
rect 313188 279822 313240 279828
rect 311912 277366 312400 277394
rect 310612 7064 310664 7070
rect 310612 7006 310664 7012
rect 311912 6730 311940 277366
rect 311900 6724 311952 6730
rect 311900 6666 311952 6672
rect 309140 6656 309192 6662
rect 309140 6598 309192 6604
rect 307760 6588 307812 6594
rect 307760 6530 307812 6536
rect 307944 6180 307996 6186
rect 307944 6122 307996 6128
rect 307024 3324 307076 3330
rect 307024 3266 307076 3272
rect 307956 480 307984 6122
rect 310244 4616 310296 4622
rect 310244 4558 310296 4564
rect 309048 3324 309100 3330
rect 309048 3266 309100 3272
rect 309060 480 309088 3266
rect 310256 480 310284 4558
rect 313200 3398 313228 279822
rect 313924 279200 313976 279206
rect 313924 279142 313976 279148
rect 313832 4480 313884 4486
rect 313832 4422 313884 4428
rect 312636 3392 312688 3398
rect 312636 3334 312688 3340
rect 313188 3392 313240 3398
rect 313188 3334 313240 3340
rect 311440 3120 311492 3126
rect 311440 3062 311492 3068
rect 311452 480 311480 3062
rect 312648 480 312676 3334
rect 313844 480 313872 4422
rect 313936 4146 313964 279142
rect 314016 278520 314068 278526
rect 314016 278462 314068 278468
rect 313924 4140 313976 4146
rect 313924 4082 313976 4088
rect 314028 3058 314056 278462
rect 314672 277642 314700 281846
rect 314660 277636 314712 277642
rect 314660 277578 314712 277584
rect 314948 277394 314976 281846
rect 316040 279336 316092 279342
rect 316040 279278 316092 279284
rect 314672 277366 314976 277394
rect 314672 6798 314700 277366
rect 316052 163606 316080 279278
rect 316144 276690 316172 281846
rect 316972 279342 317000 281846
rect 316960 279336 317012 279342
rect 316960 279278 317012 279284
rect 316684 277976 316736 277982
rect 316684 277918 316736 277924
rect 316132 276684 316184 276690
rect 316132 276626 316184 276632
rect 316040 163600 316092 163606
rect 316040 163542 316092 163548
rect 314660 6792 314712 6798
rect 314660 6734 314712 6740
rect 316224 4140 316276 4146
rect 316224 4082 316276 4088
rect 314016 3052 314068 3058
rect 314016 2994 314068 3000
rect 315028 3052 315080 3058
rect 315028 2994 315080 3000
rect 315040 480 315068 2994
rect 316236 480 316264 4082
rect 316696 2990 316724 277918
rect 317432 6866 317460 281846
rect 318812 279954 318840 281846
rect 318800 279948 318852 279954
rect 318800 279890 318852 279896
rect 317512 279608 317564 279614
rect 317512 279550 317564 279556
rect 317524 276894 317552 279550
rect 319548 277506 319576 281846
rect 320088 280152 320140 280158
rect 320088 280094 320140 280100
rect 319536 277500 319588 277506
rect 319536 277442 319588 277448
rect 317512 276888 317564 276894
rect 317512 276830 317564 276836
rect 318064 276684 318116 276690
rect 318064 276626 318116 276632
rect 317420 6860 317472 6866
rect 317420 6802 317472 6808
rect 317328 4548 317380 4554
rect 317328 4490 317380 4496
rect 316684 2984 316736 2990
rect 316684 2926 316736 2932
rect 317340 480 317368 4490
rect 318076 3058 318104 276626
rect 318524 6248 318576 6254
rect 318524 6190 318576 6196
rect 318064 3052 318116 3058
rect 318064 2994 318116 3000
rect 318536 480 318564 6190
rect 319732 598 319944 626
rect 319732 480 319760 598
rect 319916 490 319944 598
rect 320100 490 320128 280094
rect 320192 8702 320220 281846
rect 321618 281602 321646 281860
rect 321572 281574 321646 281602
rect 321756 281846 322460 281874
rect 323044 281846 323288 281874
rect 323872 281846 324208 281874
rect 324332 281846 325036 281874
rect 321572 279614 321600 281574
rect 321560 279608 321612 279614
rect 321560 279550 321612 279556
rect 320824 279132 320876 279138
rect 320824 279074 320876 279080
rect 320180 8696 320232 8702
rect 320180 8638 320232 8644
rect 320836 3194 320864 279074
rect 321756 11966 321784 281846
rect 322204 279948 322256 279954
rect 322204 279890 322256 279896
rect 321744 11960 321796 11966
rect 321744 11902 321796 11908
rect 322216 6914 322244 279890
rect 323044 11898 323072 281846
rect 323872 280022 323900 281846
rect 323860 280016 323912 280022
rect 323860 279958 323912 279964
rect 323584 279336 323636 279342
rect 323584 279278 323636 279284
rect 323032 11892 323084 11898
rect 323032 11834 323084 11840
rect 322032 6886 322244 6914
rect 320916 4412 320968 4418
rect 320916 4354 320968 4360
rect 320824 3188 320876 3194
rect 320824 3130 320876 3136
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 319916 462 320128 490
rect 320928 480 320956 4354
rect 322032 3602 322060 6886
rect 322020 3596 322072 3602
rect 322020 3538 322072 3544
rect 322112 3596 322164 3602
rect 322112 3538 322164 3544
rect 322124 480 322152 3538
rect 323308 3392 323360 3398
rect 323308 3334 323360 3340
rect 323320 480 323348 3334
rect 323596 3262 323624 279278
rect 324332 12102 324360 281846
rect 325850 281602 325878 281860
rect 326356 281846 326692 281874
rect 327184 281846 327612 281874
rect 328104 281846 328440 281874
rect 328932 281846 329268 281874
rect 329852 281846 330096 281874
rect 330680 281846 331016 281874
rect 331508 281846 331844 281874
rect 325850 281574 325924 281602
rect 325620 280126 325832 280154
rect 324964 276888 325016 276894
rect 324964 276830 325016 276836
rect 324320 12096 324372 12102
rect 324320 12038 324372 12044
rect 324412 4276 324464 4282
rect 324412 4218 324464 4224
rect 323584 3256 323636 3262
rect 323584 3198 323636 3204
rect 324424 480 324452 4218
rect 324976 3602 325004 276830
rect 325620 276758 325648 280126
rect 325804 280022 325832 280126
rect 325792 280016 325844 280022
rect 325792 279958 325844 279964
rect 325896 278050 325924 281574
rect 326356 280022 326384 281846
rect 326344 280016 326396 280022
rect 326344 279958 326396 279964
rect 327080 279608 327132 279614
rect 327080 279550 327132 279556
rect 325884 278044 325936 278050
rect 325884 277986 325936 277992
rect 325608 276752 325660 276758
rect 325608 276694 325660 276700
rect 327092 8770 327120 279550
rect 327184 12034 327212 281846
rect 328104 279614 328132 281846
rect 328932 280022 328960 281846
rect 328920 280016 328972 280022
rect 328920 279958 328972 279964
rect 329104 280016 329156 280022
rect 329104 279958 329156 279964
rect 328092 279608 328144 279614
rect 328092 279550 328144 279556
rect 327172 12028 327224 12034
rect 327172 11970 327224 11976
rect 327080 8764 327132 8770
rect 327080 8706 327132 8712
rect 328000 4344 328052 4350
rect 328000 4286 328052 4292
rect 324964 3596 325016 3602
rect 324964 3538 325016 3544
rect 326804 3460 326856 3466
rect 326804 3402 326856 3408
rect 325608 3188 325660 3194
rect 325608 3130 325660 3136
rect 325620 480 325648 3130
rect 326816 480 326844 3402
rect 328012 480 328040 4286
rect 329116 3466 329144 279958
rect 329852 278118 329880 281846
rect 329840 278112 329892 278118
rect 329840 278054 329892 278060
rect 330680 277394 330708 281846
rect 331508 279206 331536 281846
rect 332658 281602 332686 281860
rect 332612 281574 332686 281602
rect 333164 281846 333500 281874
rect 334176 281846 334420 281874
rect 334912 281846 335248 281874
rect 335372 281846 336076 281874
rect 336752 281846 336904 281874
rect 337028 281846 337824 281874
rect 338224 281846 338652 281874
rect 339052 281846 339480 281874
rect 339604 281846 340400 281874
rect 340984 281846 341228 281874
rect 341720 281846 342056 281874
rect 342272 281846 342884 281874
rect 343652 281846 343804 281874
rect 344296 281846 344632 281874
rect 345032 281846 345460 281874
rect 345676 281846 346288 281874
rect 346872 281846 347208 281874
rect 347792 281846 348036 281874
rect 348528 281846 348864 281874
rect 349172 281846 349692 281874
rect 331496 279200 331548 279206
rect 331496 279142 331548 279148
rect 332612 278254 332640 281574
rect 332600 278248 332652 278254
rect 332600 278190 332652 278196
rect 333164 278186 333192 281846
rect 334072 279608 334124 279614
rect 334072 279550 334124 279556
rect 333888 279200 333940 279206
rect 333888 279142 333940 279148
rect 333152 278180 333204 278186
rect 333152 278122 333204 278128
rect 331864 278112 331916 278118
rect 331864 278054 331916 278060
rect 329852 277366 330708 277394
rect 329852 243574 329880 277366
rect 329840 243568 329892 243574
rect 329840 243510 329892 243516
rect 329104 3460 329156 3466
rect 329104 3402 329156 3408
rect 331588 3460 331640 3466
rect 331588 3402 331640 3408
rect 329196 3392 329248 3398
rect 329196 3334 329248 3340
rect 329208 480 329236 3334
rect 330392 3256 330444 3262
rect 330392 3198 330444 3204
rect 330404 480 330432 3198
rect 331600 480 331628 3402
rect 331876 3398 331904 278054
rect 332508 278044 332560 278050
rect 332508 277986 332560 277992
rect 332520 3466 332548 277986
rect 332508 3460 332560 3466
rect 332508 3402 332560 3408
rect 331864 3392 331916 3398
rect 331864 3334 331916 3340
rect 332692 2984 332744 2990
rect 332692 2926 332744 2932
rect 332704 480 332732 2926
rect 333900 480 333928 279142
rect 334084 8974 334112 279550
rect 334072 8968 334124 8974
rect 334072 8910 334124 8916
rect 334176 3126 334204 281846
rect 334912 279614 334940 281846
rect 334900 279608 334952 279614
rect 334900 279550 334952 279556
rect 335372 9246 335400 281846
rect 336752 279478 336780 281846
rect 336740 279472 336792 279478
rect 336740 279414 336792 279420
rect 336004 277908 336056 277914
rect 336004 277850 336056 277856
rect 335360 9240 335412 9246
rect 335360 9182 335412 9188
rect 335084 6316 335136 6322
rect 335084 6258 335136 6264
rect 334164 3120 334216 3126
rect 334164 3062 334216 3068
rect 335096 480 335124 6258
rect 336016 3058 336044 277850
rect 337028 4826 337056 281846
rect 338224 277166 338252 281846
rect 339052 277394 339080 281846
rect 339408 278180 339460 278186
rect 339408 278122 339460 278128
rect 338316 277366 339080 277394
rect 338212 277160 338264 277166
rect 338212 277102 338264 277108
rect 337016 4820 337068 4826
rect 337016 4762 337068 4768
rect 338316 3534 338344 277366
rect 339420 3534 339448 278122
rect 339604 4894 339632 281846
rect 340984 277302 341012 281846
rect 341720 279546 341748 281846
rect 341708 279540 341760 279546
rect 341708 279482 341760 279488
rect 342168 279472 342220 279478
rect 342168 279414 342220 279420
rect 342076 278248 342128 278254
rect 342076 278190 342128 278196
rect 340972 277296 341024 277302
rect 340972 277238 341024 277244
rect 340144 276752 340196 276758
rect 340144 276694 340196 276700
rect 339868 6384 339920 6390
rect 339868 6326 339920 6332
rect 339592 4888 339644 4894
rect 339592 4830 339644 4836
rect 338304 3528 338356 3534
rect 338304 3470 338356 3476
rect 338672 3528 338724 3534
rect 338672 3470 338724 3476
rect 339408 3528 339460 3534
rect 339408 3470 339460 3476
rect 337476 3460 337528 3466
rect 337476 3402 337528 3408
rect 336004 3052 336056 3058
rect 336004 2994 336056 3000
rect 336280 3052 336332 3058
rect 336280 2994 336332 3000
rect 336292 480 336320 2994
rect 337488 480 337516 3402
rect 338684 480 338712 3470
rect 339880 480 339908 6326
rect 340156 3194 340184 276694
rect 342088 11898 342116 278190
rect 342076 11892 342128 11898
rect 342076 11834 342128 11840
rect 342180 11778 342208 279414
rect 341996 11750 342208 11778
rect 341996 3534 342024 11750
rect 342168 11688 342220 11694
rect 342168 11630 342220 11636
rect 340972 3528 341024 3534
rect 340972 3470 341024 3476
rect 341984 3528 342036 3534
rect 341984 3470 342036 3476
rect 340144 3188 340196 3194
rect 340144 3130 340196 3136
rect 340984 480 341012 3470
rect 342180 480 342208 11630
rect 342272 9110 342300 281846
rect 342904 279540 342956 279546
rect 342904 279482 342956 279488
rect 342260 9104 342312 9110
rect 342260 9046 342312 9052
rect 342916 3670 342944 279482
rect 343652 278390 343680 281846
rect 344296 279546 344324 281846
rect 344284 279540 344336 279546
rect 344284 279482 344336 279488
rect 343640 278384 343692 278390
rect 343640 278326 343692 278332
rect 343364 7812 343416 7818
rect 343364 7754 343416 7760
rect 342904 3664 342956 3670
rect 342904 3606 342956 3612
rect 343376 480 343404 7754
rect 345032 4962 345060 281846
rect 345676 277394 345704 281846
rect 346872 279342 346900 281846
rect 346860 279336 346912 279342
rect 346860 279278 346912 279284
rect 345124 277366 345704 277394
rect 345124 9178 345152 277366
rect 347044 277160 347096 277166
rect 347044 277102 347096 277108
rect 345112 9172 345164 9178
rect 345112 9114 345164 9120
rect 347056 6914 347084 277102
rect 346872 6886 347084 6914
rect 345756 6452 345808 6458
rect 345756 6394 345808 6400
rect 345020 4956 345072 4962
rect 345020 4898 345072 4904
rect 344560 3188 344612 3194
rect 344560 3130 344612 3136
rect 344572 480 344600 3130
rect 345768 480 345796 6394
rect 346872 2990 346900 6886
rect 347792 5098 347820 281846
rect 348528 278322 348556 281846
rect 349068 279540 349120 279546
rect 349068 279482 349120 279488
rect 348516 278316 348568 278322
rect 348516 278258 348568 278264
rect 347780 5092 347832 5098
rect 347780 5034 347832 5040
rect 349080 3534 349108 279482
rect 349172 3738 349200 281846
rect 350598 281602 350626 281860
rect 350552 281574 350626 281602
rect 351104 281846 351440 281874
rect 351932 281846 352268 281874
rect 352392 281846 353096 281874
rect 353312 281846 354016 281874
rect 354692 281846 354844 281874
rect 355336 281846 355672 281874
rect 356164 281846 356500 281874
rect 357084 281846 357420 281874
rect 357544 281846 358248 281874
rect 358924 281846 359076 281874
rect 359568 281846 359904 281874
rect 360212 281846 360824 281874
rect 349804 278792 349856 278798
rect 349804 278734 349856 278740
rect 349816 3942 349844 278734
rect 350448 93152 350500 93158
rect 350448 93094 350500 93100
rect 349804 3936 349856 3942
rect 349804 3878 349856 3884
rect 349160 3732 349212 3738
rect 349160 3674 349212 3680
rect 350460 3534 350488 93094
rect 350552 5030 350580 281574
rect 351104 278730 351132 281846
rect 351932 280158 351960 281846
rect 351920 280152 351972 280158
rect 351920 280094 351972 280100
rect 351092 278724 351144 278730
rect 351092 278666 351144 278672
rect 352392 277394 352420 281846
rect 352564 280152 352616 280158
rect 352564 280094 352616 280100
rect 352024 277366 352420 277394
rect 352024 9042 352052 277366
rect 352012 9036 352064 9042
rect 352012 8978 352064 8984
rect 350540 5024 350592 5030
rect 350540 4966 350592 4972
rect 351644 3664 351696 3670
rect 351644 3606 351696 3612
rect 348056 3528 348108 3534
rect 348056 3470 348108 3476
rect 349068 3528 349120 3534
rect 349068 3470 349120 3476
rect 349252 3528 349304 3534
rect 349252 3470 349304 3476
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 346860 2984 346912 2990
rect 346860 2926 346912 2932
rect 346952 2984 347004 2990
rect 346952 2926 347004 2932
rect 346964 480 346992 2926
rect 348068 480 348096 3470
rect 349264 480 349292 3470
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 350460 480 350488 3334
rect 351656 480 351684 3606
rect 352576 3398 352604 280094
rect 353312 10470 353340 281846
rect 354692 278798 354720 281846
rect 354680 278792 354732 278798
rect 354680 278734 354732 278740
rect 355336 278458 355364 281846
rect 355324 278452 355376 278458
rect 355324 278394 355376 278400
rect 353944 278316 353996 278322
rect 353944 278258 353996 278264
rect 353300 10464 353352 10470
rect 353300 10406 353352 10412
rect 353956 3942 353984 278258
rect 356164 277098 356192 281846
rect 357084 279410 357112 281846
rect 357072 279404 357124 279410
rect 357072 279346 357124 279352
rect 356704 279200 356756 279206
rect 356704 279142 356756 279148
rect 356152 277092 356204 277098
rect 356152 277034 356204 277040
rect 352840 3936 352892 3942
rect 352840 3878 352892 3884
rect 353944 3936 353996 3942
rect 353944 3878 353996 3884
rect 356336 3936 356388 3942
rect 356336 3878 356388 3884
rect 352564 3392 352616 3398
rect 352564 3334 352616 3340
rect 352852 480 352880 3878
rect 355232 3800 355284 3806
rect 355232 3742 355284 3748
rect 354036 3732 354088 3738
rect 354036 3674 354088 3680
rect 354048 480 354076 3674
rect 355244 480 355272 3742
rect 356348 480 356376 3878
rect 356716 3806 356744 279142
rect 357348 278384 357400 278390
rect 357348 278326 357400 278332
rect 357360 3942 357388 278326
rect 357544 6118 357572 281846
rect 358820 279404 358872 279410
rect 358820 279346 358872 279352
rect 358728 279336 358780 279342
rect 358728 279278 358780 279284
rect 357532 6112 357584 6118
rect 357532 6054 357584 6060
rect 358740 3942 358768 279278
rect 357348 3936 357400 3942
rect 357348 3878 357400 3884
rect 357532 3936 357584 3942
rect 357532 3878 357584 3884
rect 358728 3936 358780 3942
rect 358728 3878 358780 3884
rect 356704 3800 356756 3806
rect 356704 3742 356756 3748
rect 357544 480 357572 3878
rect 358636 3868 358688 3874
rect 358636 3810 358688 3816
rect 358648 1986 358676 3810
rect 358832 3398 358860 279346
rect 358924 276826 358952 281846
rect 359568 279410 359596 281846
rect 359556 279404 359608 279410
rect 359556 279346 359608 279352
rect 360108 278452 360160 278458
rect 360108 278394 360160 278400
rect 358912 276820 358964 276826
rect 358912 276762 358964 276768
rect 358820 3392 358872 3398
rect 358820 3334 358872 3340
rect 360120 2774 360148 278394
rect 360212 6050 360240 281846
rect 361638 281602 361666 281860
rect 361592 281574 361666 281602
rect 362144 281846 362480 281874
rect 362972 281846 363400 281874
rect 363524 281846 364228 281874
rect 364720 281846 365056 281874
rect 365732 281846 365884 281874
rect 366468 281846 366804 281874
rect 367296 281846 367632 281874
rect 367756 281846 368460 281874
rect 368952 281846 369288 281874
rect 369872 281846 370208 281874
rect 370332 281846 371036 281874
rect 371252 281846 371864 281874
rect 361592 277030 361620 281574
rect 362144 279274 362172 281846
rect 362132 279268 362184 279274
rect 362132 279210 362184 279216
rect 361580 277024 361632 277030
rect 361580 276966 361632 276972
rect 360844 276820 360896 276826
rect 360844 276762 360896 276768
rect 360200 6044 360252 6050
rect 360200 5986 360252 5992
rect 360856 3058 360884 276762
rect 362972 5982 363000 281846
rect 363524 277394 363552 281846
rect 364720 278798 364748 281846
rect 364984 279268 365036 279274
rect 364984 279210 365036 279216
rect 363604 278792 363656 278798
rect 363604 278734 363656 278740
rect 364708 278792 364760 278798
rect 364708 278734 364760 278740
rect 363064 277366 363552 277394
rect 363064 276962 363092 277366
rect 363052 276956 363104 276962
rect 363052 276898 363104 276904
rect 362960 5976 363012 5982
rect 362960 5918 363012 5924
rect 363616 3806 363644 278734
rect 364248 278724 364300 278730
rect 364248 278666 364300 278672
rect 363604 3800 363656 3806
rect 363604 3742 363656 3748
rect 364260 3398 364288 278666
rect 363512 3392 363564 3398
rect 363512 3334 363564 3340
rect 364248 3392 364300 3398
rect 364248 3334 364300 3340
rect 364616 3392 364668 3398
rect 364616 3334 364668 3340
rect 361120 3120 361172 3126
rect 361120 3062 361172 3068
rect 360844 3052 360896 3058
rect 360844 2994 360896 3000
rect 359936 2746 360148 2774
rect 358648 1958 358768 1986
rect 358740 480 358768 1958
rect 359936 480 359964 2746
rect 361132 480 361160 3062
rect 362316 3052 362368 3058
rect 362316 2994 362368 3000
rect 362328 480 362356 2994
rect 363524 480 363552 3334
rect 364628 480 364656 3334
rect 364996 3058 365024 279210
rect 365732 5234 365760 281846
rect 366364 279200 366416 279206
rect 366364 279142 366416 279148
rect 365720 5228 365772 5234
rect 365720 5170 365772 5176
rect 366376 3398 366404 279142
rect 366468 278662 366496 281846
rect 367296 280090 367324 281846
rect 367284 280084 367336 280090
rect 367284 280026 367336 280032
rect 367756 279698 367784 281846
rect 367204 279670 367784 279698
rect 366456 278656 366508 278662
rect 366456 278598 366508 278604
rect 367204 5302 367232 279670
rect 367744 278656 367796 278662
rect 367744 278598 367796 278604
rect 367192 5296 367244 5302
rect 367192 5238 367244 5244
rect 367756 3398 367784 278598
rect 368952 278594 368980 281846
rect 369768 280084 369820 280090
rect 369768 280026 369820 280032
rect 368940 278588 368992 278594
rect 368940 278530 368992 278536
rect 368204 3800 368256 3806
rect 368204 3742 368256 3748
rect 366364 3392 366416 3398
rect 366364 3334 366416 3340
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367744 3392 367796 3398
rect 367744 3334 367796 3340
rect 364984 3052 365036 3058
rect 364984 2994 365036 3000
rect 365812 3052 365864 3058
rect 365812 2994 365864 3000
rect 365824 480 365852 2994
rect 367020 480 367048 3334
rect 368216 480 368244 3742
rect 369412 598 369624 626
rect 369412 480 369440 598
rect 369596 490 369624 598
rect 369780 490 369808 280026
rect 369872 4010 369900 281846
rect 370332 277394 370360 281846
rect 369964 277366 370360 277394
rect 369964 5370 369992 277366
rect 371252 7614 371280 281846
rect 372678 281602 372706 281860
rect 372632 281574 372706 281602
rect 372816 281846 373612 281874
rect 374104 281846 374440 281874
rect 374564 281846 375268 281874
rect 375392 281846 376096 281874
rect 376864 281846 377016 281874
rect 377508 281846 377844 281874
rect 378152 281846 378672 281874
rect 379164 281846 379500 281874
rect 379716 281846 380420 281874
rect 380912 281846 381248 281874
rect 381464 281846 382076 281874
rect 382568 281846 382904 281874
rect 372632 279682 372660 281574
rect 372620 279676 372672 279682
rect 372620 279618 372672 279624
rect 371240 7608 371292 7614
rect 371240 7550 371292 7556
rect 372816 5438 372844 281846
rect 373264 279676 373316 279682
rect 373264 279618 373316 279624
rect 372804 5432 372856 5438
rect 372804 5374 372856 5380
rect 369952 5364 370004 5370
rect 369952 5306 370004 5312
rect 370596 4820 370648 4826
rect 370596 4762 370648 4768
rect 369860 4004 369912 4010
rect 369860 3946 369912 3952
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 369596 462 369808 490
rect 370608 480 370636 4762
rect 373276 3398 373304 279618
rect 374104 277982 374132 281846
rect 374092 277976 374144 277982
rect 374092 277918 374144 277924
rect 374564 277394 374592 281846
rect 375288 278588 375340 278594
rect 375288 278530 375340 278536
rect 374012 277366 374592 277394
rect 374012 4078 374040 277366
rect 374000 4072 374052 4078
rect 374000 4014 374052 4020
rect 375196 3868 375248 3874
rect 375196 3810 375248 3816
rect 371700 3392 371752 3398
rect 371700 3334 371752 3340
rect 373264 3392 373316 3398
rect 373264 3334 373316 3340
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 371712 480 371740 3334
rect 372896 2984 372948 2990
rect 372896 2926 372948 2932
rect 372908 480 372936 2926
rect 374104 480 374132 3334
rect 375208 1986 375236 3810
rect 375300 3398 375328 278530
rect 375392 5166 375420 281846
rect 376864 7682 376892 281846
rect 377508 279750 377536 281846
rect 377496 279744 377548 279750
rect 377496 279686 377548 279692
rect 377588 279744 377640 279750
rect 377588 279686 377640 279692
rect 377600 277394 377628 279686
rect 377416 277366 377628 277394
rect 376852 7676 376904 7682
rect 376852 7618 376904 7624
rect 375380 5160 375432 5166
rect 375380 5102 375432 5108
rect 377416 3398 377444 277366
rect 377680 7608 377732 7614
rect 377680 7550 377732 7556
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 376484 3392 376536 3398
rect 376484 3334 376536 3340
rect 377404 3392 377456 3398
rect 377404 3334 377456 3340
rect 375208 1958 375328 1986
rect 375300 480 375328 1958
rect 376496 480 376524 3334
rect 377692 480 377720 7550
rect 378152 4758 378180 281846
rect 379164 278526 379192 281846
rect 379428 279132 379480 279138
rect 379428 279074 379480 279080
rect 379152 278520 379204 278526
rect 379152 278462 379204 278468
rect 378140 4752 378192 4758
rect 378140 4694 378192 4700
rect 379440 3398 379468 279074
rect 378876 3392 378928 3398
rect 378876 3334 378928 3340
rect 379428 3392 379480 3398
rect 379428 3334 379480 3340
rect 378888 480 378916 3334
rect 379716 2922 379744 281846
rect 380912 5506 380940 281846
rect 381464 277394 381492 281846
rect 382568 279818 382596 281846
rect 383810 281602 383838 281860
rect 383764 281574 383838 281602
rect 384316 281846 384652 281874
rect 385052 281846 385480 281874
rect 385788 281846 386400 281874
rect 386892 281846 387228 281874
rect 387812 281846 388056 281874
rect 388272 281846 388884 281874
rect 389192 281846 389804 281874
rect 382556 279812 382608 279818
rect 382556 279754 382608 279760
rect 383016 278792 383068 278798
rect 383016 278734 383068 278740
rect 382924 278520 382976 278526
rect 382924 278462 382976 278468
rect 381004 277366 381492 277394
rect 381004 7750 381032 277366
rect 380992 7744 381044 7750
rect 380992 7686 381044 7692
rect 380900 5500 380952 5506
rect 380900 5442 380952 5448
rect 382372 4004 382424 4010
rect 382372 3946 382424 3952
rect 381176 3392 381228 3398
rect 381176 3334 381228 3340
rect 379704 2916 379756 2922
rect 379704 2858 379756 2864
rect 379980 2916 380032 2922
rect 379980 2858 380032 2864
rect 379992 480 380020 2858
rect 381188 480 381216 3334
rect 382384 480 382412 3946
rect 382936 3398 382964 278462
rect 383028 6186 383056 278734
rect 383016 6180 383068 6186
rect 383016 6122 383068 6128
rect 383764 4690 383792 281574
rect 384316 278798 384344 281846
rect 384396 279812 384448 279818
rect 384396 279754 384448 279760
rect 384304 278792 384356 278798
rect 384304 278734 384356 278740
rect 384408 277394 384436 279754
rect 384316 277366 384436 277394
rect 383752 4684 383804 4690
rect 383752 4626 383804 4632
rect 384316 4078 384344 277366
rect 384764 4888 384816 4894
rect 384764 4830 384816 4836
rect 383568 4072 383620 4078
rect 383568 4014 383620 4020
rect 384304 4072 384356 4078
rect 384304 4014 384356 4020
rect 382924 3392 382976 3398
rect 382924 3334 382976 3340
rect 383580 480 383608 4014
rect 384776 480 384804 4830
rect 385052 3330 385080 281846
rect 385788 277394 385816 281846
rect 386892 277914 386920 281846
rect 387812 279886 387840 281846
rect 387800 279880 387852 279886
rect 387800 279822 387852 279828
rect 386880 277908 386932 277914
rect 386880 277850 386932 277856
rect 388272 277394 388300 281846
rect 388444 279064 388496 279070
rect 388444 279006 388496 279012
rect 385144 277366 385816 277394
rect 387904 277366 388300 277394
rect 385144 4622 385172 277366
rect 385132 4616 385184 4622
rect 385132 4558 385184 4564
rect 387904 4486 387932 277366
rect 387892 4480 387944 4486
rect 387892 4422 387944 4428
rect 388456 4078 388484 279006
rect 389192 276690 389220 281846
rect 390618 281602 390646 281860
rect 390572 281574 390646 281602
rect 390756 281846 391460 281874
rect 392044 281846 392288 281874
rect 392872 281846 393208 281874
rect 393332 281846 394036 281874
rect 390572 279818 390600 281574
rect 389824 279812 389876 279818
rect 389824 279754 389876 279760
rect 390560 279812 390612 279818
rect 390560 279754 390612 279760
rect 389180 276684 389232 276690
rect 389180 276626 389232 276632
rect 389836 4146 389864 279754
rect 389916 277908 389968 277914
rect 389916 277850 389968 277856
rect 389824 4140 389876 4146
rect 389824 4082 389876 4088
rect 385960 4072 386012 4078
rect 385960 4014 386012 4020
rect 388444 4072 388496 4078
rect 388444 4014 388496 4020
rect 389456 4072 389508 4078
rect 389456 4014 389508 4020
rect 385040 3324 385092 3330
rect 385040 3266 385092 3272
rect 385972 480 386000 4014
rect 388260 3324 388312 3330
rect 388260 3266 388312 3272
rect 387156 2916 387208 2922
rect 387156 2858 387208 2864
rect 387168 480 387196 2858
rect 388272 480 388300 3266
rect 389468 480 389496 4014
rect 389928 3330 389956 277850
rect 390756 4554 390784 281846
rect 391848 278996 391900 279002
rect 391848 278938 391900 278944
rect 391860 6914 391888 278938
rect 391768 6886 391888 6914
rect 390744 4548 390796 4554
rect 390744 4490 390796 4496
rect 391768 3330 391796 6886
rect 392044 6254 392072 281846
rect 392872 279954 392900 281846
rect 392860 279948 392912 279954
rect 392860 279890 392912 279896
rect 392584 277976 392636 277982
rect 392584 277918 392636 277924
rect 392032 6248 392084 6254
rect 392032 6190 392084 6196
rect 392596 3330 392624 277918
rect 393332 4418 393360 281846
rect 394850 281602 394878 281860
rect 394804 281574 394878 281602
rect 395356 281846 395692 281874
rect 396092 281846 396612 281874
rect 396736 281846 397440 281874
rect 397932 281846 398268 281874
rect 398852 281846 399096 281874
rect 399680 281846 400016 281874
rect 400232 281846 400844 281874
rect 393964 279948 394016 279954
rect 393964 279890 394016 279896
rect 393320 4412 393372 4418
rect 393320 4354 393372 4360
rect 393976 4146 394004 279890
rect 394700 279880 394752 279886
rect 394700 279822 394752 279828
rect 393044 4140 393096 4146
rect 393044 4082 393096 4088
rect 393964 4140 394016 4146
rect 393964 4082 394016 4088
rect 389916 3324 389968 3330
rect 389916 3266 389968 3272
rect 390652 3324 390704 3330
rect 390652 3266 390704 3272
rect 391756 3324 391808 3330
rect 391756 3266 391808 3272
rect 391848 3324 391900 3330
rect 391848 3266 391900 3272
rect 392584 3324 392636 3330
rect 392584 3266 392636 3272
rect 390664 480 390692 3266
rect 391860 480 391888 3266
rect 393056 480 393084 4082
rect 394712 3602 394740 279822
rect 394804 276894 394832 281574
rect 395356 279886 395384 281846
rect 395344 279880 395396 279886
rect 395344 279822 395396 279828
rect 394792 276888 394844 276894
rect 394792 276830 394844 276836
rect 396092 4282 396120 281846
rect 396736 279596 396764 281846
rect 397932 280022 397960 281846
rect 397920 280016 397972 280022
rect 397920 279958 397972 279964
rect 396184 279568 396764 279596
rect 396184 276758 396212 279568
rect 396724 277840 396776 277846
rect 396724 277782 396776 277788
rect 396172 276752 396224 276758
rect 396172 276694 396224 276700
rect 396080 4276 396132 4282
rect 396080 4218 396132 4224
rect 396736 3602 396764 277782
rect 398852 4350 398880 281846
rect 399484 280016 399536 280022
rect 399484 279958 399536 279964
rect 398840 4344 398892 4350
rect 398840 4286 398892 4292
rect 399496 3602 399524 279958
rect 399680 278118 399708 281846
rect 400128 279948 400180 279954
rect 400128 279890 400180 279896
rect 399668 278112 399720 278118
rect 399668 278054 399720 278060
rect 394700 3596 394752 3602
rect 394700 3538 394752 3544
rect 395344 3596 395396 3602
rect 395344 3538 395396 3544
rect 396724 3596 396776 3602
rect 396724 3538 396776 3544
rect 397736 3596 397788 3602
rect 397736 3538 397788 3544
rect 399484 3596 399536 3602
rect 399484 3538 399536 3544
rect 394240 2916 394292 2922
rect 394240 2858 394292 2864
rect 394252 480 394280 2858
rect 395356 480 395384 3538
rect 396540 2848 396592 2854
rect 396540 2790 396592 2796
rect 396552 480 396580 2790
rect 397748 480 397776 3538
rect 398932 3256 398984 3262
rect 398932 3198 398984 3204
rect 398944 480 398972 3198
rect 400140 480 400168 279890
rect 400232 4146 400260 281846
rect 401658 281602 401686 281860
rect 401612 281574 401686 281602
rect 401796 281846 402500 281874
rect 403176 281846 403420 281874
rect 403544 281846 404248 281874
rect 404372 281846 405076 281874
rect 400864 278112 400916 278118
rect 400864 278054 400916 278060
rect 400220 4140 400272 4146
rect 400220 4082 400272 4088
rect 400876 3262 400904 278054
rect 401612 278050 401640 281574
rect 401600 278044 401652 278050
rect 401600 277986 401652 277992
rect 401796 277166 401824 281846
rect 403176 279614 403204 281846
rect 403164 279608 403216 279614
rect 403164 279550 403216 279556
rect 403544 277394 403572 281846
rect 403624 278044 403676 278050
rect 403624 277986 403676 277992
rect 403084 277366 403572 277394
rect 401784 277160 401836 277166
rect 401784 277102 401836 277108
rect 403084 6322 403112 277366
rect 403636 6914 403664 277986
rect 404372 276826 404400 281846
rect 405890 281602 405918 281860
rect 405844 281574 405918 281602
rect 406488 281846 406824 281874
rect 407224 281846 407652 281874
rect 408144 281846 408480 281874
rect 409064 281846 409400 281874
rect 409984 281846 410228 281874
rect 410720 281846 411056 281874
rect 411272 281846 411884 281874
rect 405648 278860 405700 278866
rect 405648 278802 405700 278808
rect 404360 276820 404412 276826
rect 404360 276762 404412 276768
rect 403176 6886 403664 6914
rect 403072 6316 403124 6322
rect 403072 6258 403124 6264
rect 401324 4140 401376 4146
rect 401324 4082 401376 4088
rect 402520 4140 402572 4146
rect 402520 4082 402572 4088
rect 402980 4140 403032 4146
rect 403176 4128 403204 6886
rect 403032 4100 403204 4128
rect 402980 4082 403032 4088
rect 400864 3256 400916 3262
rect 400864 3198 400916 3204
rect 401336 480 401364 4082
rect 402532 480 402560 4082
rect 405660 3534 405688 278802
rect 404820 3528 404872 3534
rect 404820 3470 404872 3476
rect 405648 3528 405700 3534
rect 405648 3470 405700 3476
rect 403624 3256 403676 3262
rect 403624 3198 403676 3204
rect 403636 480 403664 3198
rect 404832 480 404860 3470
rect 405844 3466 405872 281574
rect 406488 278186 406516 281846
rect 406476 278180 406528 278186
rect 406476 278122 406528 278128
rect 407028 278180 407080 278186
rect 407028 278122 407080 278128
rect 407040 3534 407068 278122
rect 407224 6390 407252 281846
rect 407764 279608 407816 279614
rect 407764 279550 407816 279556
rect 407212 6384 407264 6390
rect 407212 6326 407264 6332
rect 406016 3528 406068 3534
rect 406016 3470 406068 3476
rect 407028 3528 407080 3534
rect 407028 3470 407080 3476
rect 407212 3528 407264 3534
rect 407212 3470 407264 3476
rect 405832 3460 405884 3466
rect 405832 3402 405884 3408
rect 406028 480 406056 3470
rect 407224 480 407252 3470
rect 407776 3194 407804 279550
rect 408144 279478 408172 281846
rect 408132 279472 408184 279478
rect 408132 279414 408184 279420
rect 409064 278254 409092 281846
rect 409144 278928 409196 278934
rect 409144 278870 409196 278876
rect 409052 278248 409104 278254
rect 409052 278190 409104 278196
rect 409156 3534 409184 278870
rect 409984 7818 410012 281846
rect 410720 279614 410748 281846
rect 410708 279608 410760 279614
rect 410708 279550 410760 279556
rect 410524 278248 410576 278254
rect 410524 278190 410576 278196
rect 409972 7812 410024 7818
rect 409972 7754 410024 7760
rect 410536 3534 410564 278190
rect 411272 6458 411300 281846
rect 412790 281602 412818 281860
rect 412744 281574 412818 281602
rect 413296 281846 413632 281874
rect 414124 281846 414460 281874
rect 414952 281846 415288 281874
rect 415412 281846 416208 281874
rect 416792 281846 417036 281874
rect 417160 281846 417864 281874
rect 418356 281846 418692 281874
rect 412548 279472 412600 279478
rect 412548 279414 412600 279420
rect 411260 6452 411312 6458
rect 411260 6394 411312 6400
rect 412560 3534 412588 279414
rect 409144 3528 409196 3534
rect 409144 3470 409196 3476
rect 409604 3528 409656 3534
rect 409604 3470 409656 3476
rect 410524 3528 410576 3534
rect 410524 3470 410576 3476
rect 411904 3528 411956 3534
rect 411904 3470 411956 3476
rect 412548 3528 412600 3534
rect 412548 3470 412600 3476
rect 408408 3460 408460 3466
rect 408408 3402 408460 3408
rect 407764 3188 407816 3194
rect 407764 3130 407816 3136
rect 408420 480 408448 3402
rect 409616 480 409644 3470
rect 410800 3188 410852 3194
rect 410800 3130 410852 3136
rect 410812 480 410840 3130
rect 411916 480 411944 3470
rect 412744 2854 412772 281574
rect 413296 279546 413324 281846
rect 413284 279540 413336 279546
rect 413284 279482 413336 279488
rect 413928 277772 413980 277778
rect 413928 277714 413980 277720
rect 413940 3534 413968 277714
rect 414124 93158 414152 281846
rect 414952 280158 414980 281846
rect 414940 280152 414992 280158
rect 414940 280094 414992 280100
rect 415308 279540 415360 279546
rect 415308 279482 415360 279488
rect 414112 93152 414164 93158
rect 414112 93094 414164 93100
rect 415320 3534 415348 279482
rect 415412 3670 415440 281846
rect 416792 278322 416820 281846
rect 416780 278316 416832 278322
rect 416780 278258 416832 278264
rect 417160 277394 417188 281846
rect 418356 279410 418384 281846
rect 419598 281602 419626 281860
rect 419552 281574 419626 281602
rect 420104 281846 420440 281874
rect 420932 281846 421268 281874
rect 421760 281846 422096 281874
rect 422680 281846 423016 281874
rect 423692 281846 423844 281874
rect 424244 281846 424672 281874
rect 425164 281846 425500 281874
rect 426084 281846 426420 281874
rect 426912 281846 427248 281874
rect 427924 281846 428076 281874
rect 428660 281846 428996 281874
rect 429212 281846 429824 281874
rect 419448 280152 419500 280158
rect 419448 280094 419500 280100
rect 418344 279404 418396 279410
rect 418344 279346 418396 279352
rect 417424 278316 417476 278322
rect 417424 278258 417476 278264
rect 416792 277366 417188 277394
rect 416792 3738 416820 277366
rect 416780 3732 416832 3738
rect 416780 3674 416832 3680
rect 415400 3664 415452 3670
rect 415400 3606 415452 3612
rect 417436 3534 417464 278258
rect 419460 3534 419488 280094
rect 419552 278390 419580 281574
rect 420104 279342 420132 281846
rect 420092 279336 420144 279342
rect 420092 279278 420144 279284
rect 420184 278792 420236 278798
rect 420184 278734 420236 278740
rect 419540 278384 419592 278390
rect 419540 278326 419592 278332
rect 420196 6914 420224 278734
rect 420104 6886 420224 6914
rect 413100 3528 413152 3534
rect 413100 3470 413152 3476
rect 413928 3528 413980 3534
rect 413928 3470 413980 3476
rect 414296 3528 414348 3534
rect 414296 3470 414348 3476
rect 415308 3528 415360 3534
rect 415308 3470 415360 3476
rect 416688 3528 416740 3534
rect 416688 3470 416740 3476
rect 417424 3528 417476 3534
rect 417424 3470 417476 3476
rect 418988 3528 419040 3534
rect 418988 3470 419040 3476
rect 419448 3528 419500 3534
rect 419448 3470 419500 3476
rect 412732 2848 412784 2854
rect 412732 2790 412784 2796
rect 413112 480 413140 3470
rect 414308 480 414336 3470
rect 415492 3120 415544 3126
rect 415492 3062 415544 3068
rect 415504 480 415532 3062
rect 416700 480 416728 3470
rect 417884 2848 417936 2854
rect 417884 2790 417936 2796
rect 417896 480 417924 2790
rect 419000 480 419028 3470
rect 420104 3058 420132 6886
rect 420932 3942 420960 281846
rect 421564 279404 421616 279410
rect 421564 279346 421616 279352
rect 420920 3936 420972 3942
rect 420920 3878 420972 3884
rect 420184 3732 420236 3738
rect 420184 3674 420236 3680
rect 421380 3732 421432 3738
rect 421380 3674 421432 3680
rect 420092 3052 420144 3058
rect 420092 2994 420144 3000
rect 420196 480 420224 3674
rect 421392 480 421420 3674
rect 421576 3670 421604 279346
rect 421760 278458 421788 281846
rect 422680 278798 422708 281846
rect 423692 279274 423720 281846
rect 423680 279268 423732 279274
rect 423680 279210 423732 279216
rect 422668 278792 422720 278798
rect 422668 278734 422720 278740
rect 424244 278730 424272 281846
rect 425164 279206 425192 281846
rect 425704 279676 425756 279682
rect 425704 279618 425756 279624
rect 425152 279200 425204 279206
rect 425152 279142 425204 279148
rect 424232 278724 424284 278730
rect 424232 278666 424284 278672
rect 424324 278724 424376 278730
rect 424324 278666 424376 278672
rect 421748 278452 421800 278458
rect 421748 278394 421800 278400
rect 424336 3942 424364 278666
rect 424324 3936 424376 3942
rect 424324 3878 424376 3884
rect 421564 3664 421616 3670
rect 421564 3606 421616 3612
rect 424968 3664 425020 3670
rect 424968 3606 425020 3612
rect 423772 3392 423824 3398
rect 423772 3334 423824 3340
rect 422576 3120 422628 3126
rect 422576 3062 422628 3068
rect 422588 480 422616 3062
rect 423784 480 423812 3334
rect 424980 480 425008 3606
rect 425716 2990 425744 279618
rect 426084 279410 426112 281846
rect 426072 279404 426124 279410
rect 426072 279346 426124 279352
rect 426912 278662 426940 281846
rect 426900 278656 426952 278662
rect 426900 278598 426952 278604
rect 425796 278452 425848 278458
rect 425796 278394 425848 278400
rect 425808 3398 425836 278394
rect 427924 3806 427952 281846
rect 428660 280090 428688 281846
rect 428648 280084 428700 280090
rect 428648 280026 428700 280032
rect 428464 278384 428516 278390
rect 428464 278326 428516 278332
rect 427912 3800 427964 3806
rect 427912 3742 427964 3748
rect 428476 3398 428504 278326
rect 429212 4826 429240 281846
rect 430638 281602 430666 281860
rect 430592 281574 430666 281602
rect 431144 281846 431480 281874
rect 432064 281846 432400 281874
rect 432616 281846 433228 281874
rect 433720 281846 434056 281874
rect 430488 280084 430540 280090
rect 430488 280026 430540 280032
rect 429200 4820 429252 4826
rect 429200 4762 429252 4768
rect 430500 3398 430528 280026
rect 430592 279342 430620 281574
rect 431144 279682 431172 281846
rect 431132 279676 431184 279682
rect 431132 279618 431184 279624
rect 431224 279404 431276 279410
rect 431224 279346 431276 279352
rect 430580 279336 430632 279342
rect 430580 279278 430632 279284
rect 431236 3942 431264 279346
rect 432064 278594 432092 281846
rect 432052 278588 432104 278594
rect 432052 278530 432104 278536
rect 432616 277394 432644 281846
rect 433720 279750 433748 281846
rect 434870 281602 434898 281860
rect 434824 281574 434898 281602
rect 435468 281846 435804 281874
rect 436296 281846 436632 281874
rect 437124 281846 437460 281874
rect 437676 281846 438288 281874
rect 438872 281846 439208 281874
rect 439608 281846 440036 281874
rect 440528 281846 440864 281874
rect 433708 279744 433760 279750
rect 433708 279686 433760 279692
rect 433248 279676 433300 279682
rect 433248 279618 433300 279624
rect 431972 277366 432644 277394
rect 431868 276684 431920 276690
rect 431868 276626 431920 276632
rect 431224 3936 431276 3942
rect 431224 3878 431276 3884
rect 431880 3398 431908 276626
rect 431972 3874 432000 277366
rect 431960 3868 432012 3874
rect 431960 3810 432012 3816
rect 433260 3398 433288 279618
rect 434824 7614 434852 281574
rect 435468 279138 435496 281846
rect 436296 279410 436324 281846
rect 436284 279404 436336 279410
rect 436284 279346 436336 279352
rect 435456 279132 435508 279138
rect 435456 279074 435508 279080
rect 436744 278792 436796 278798
rect 436744 278734 436796 278740
rect 435364 278588 435416 278594
rect 435364 278530 435416 278536
rect 434812 7608 434864 7614
rect 434812 7550 434864 7556
rect 425796 3392 425848 3398
rect 425796 3334 425848 3340
rect 427268 3392 427320 3398
rect 427268 3334 427320 3340
rect 428464 3392 428516 3398
rect 428464 3334 428516 3340
rect 429660 3392 429712 3398
rect 429660 3334 429712 3340
rect 430488 3392 430540 3398
rect 430488 3334 430540 3340
rect 430856 3392 430908 3398
rect 430856 3334 430908 3340
rect 431868 3392 431920 3398
rect 431868 3334 431920 3340
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 425704 2984 425756 2990
rect 425704 2926 425756 2932
rect 426164 2984 426216 2990
rect 426164 2926 426216 2932
rect 426176 480 426204 2926
rect 427280 480 427308 3334
rect 428464 3052 428516 3058
rect 428464 2994 428516 3000
rect 428476 480 428504 2994
rect 429672 480 429700 3334
rect 430868 480 430896 3334
rect 432064 480 432092 3334
rect 435376 3330 435404 278530
rect 436756 6914 436784 278734
rect 437124 278526 437152 281846
rect 437388 279744 437440 279750
rect 437388 279686 437440 279692
rect 437112 278520 437164 278526
rect 437112 278462 437164 278468
rect 436664 6886 436784 6914
rect 436664 3398 436692 6886
rect 437400 3398 437428 279686
rect 437676 4010 437704 281846
rect 438872 279818 438900 281846
rect 438860 279812 438912 279818
rect 438860 279754 438912 279760
rect 439608 277394 439636 281846
rect 440148 279812 440200 279818
rect 440148 279754 440200 279760
rect 438964 277366 439636 277394
rect 438964 4894 438992 277366
rect 438952 4888 439004 4894
rect 438952 4830 439004 4836
rect 437664 4004 437716 4010
rect 437664 3946 437716 3952
rect 440160 3398 440188 279754
rect 440528 279070 440556 281846
rect 441678 281602 441706 281860
rect 441632 281574 441706 281602
rect 442368 281846 442612 281874
rect 443104 281846 443440 281874
rect 443932 281846 444268 281874
rect 444760 281846 445096 281874
rect 445772 281846 446016 281874
rect 446508 281846 446844 281874
rect 447336 281846 447672 281874
rect 447796 281846 448500 281874
rect 449084 281846 449420 281874
rect 449912 281846 450248 281874
rect 450740 281846 451076 281874
rect 451292 281846 451996 281874
rect 452672 281846 452824 281874
rect 452948 281846 453652 281874
rect 454144 281846 454480 281874
rect 455064 281846 455400 281874
rect 455892 281846 456228 281874
rect 440516 279064 440568 279070
rect 440516 279006 440568 279012
rect 441632 278798 441660 281574
rect 442264 278996 442316 279002
rect 442264 278938 442316 278944
rect 441620 278792 441672 278798
rect 441620 278734 441672 278740
rect 440884 278520 440936 278526
rect 440884 278462 440936 278468
rect 440332 4004 440384 4010
rect 440332 3946 440384 3952
rect 436652 3392 436704 3398
rect 436652 3334 436704 3340
rect 436744 3392 436796 3398
rect 436744 3334 436796 3340
rect 437388 3392 437440 3398
rect 437388 3334 437440 3340
rect 439136 3392 439188 3398
rect 439136 3334 439188 3340
rect 440148 3392 440200 3398
rect 440148 3334 440200 3340
rect 434444 3324 434496 3330
rect 434444 3266 434496 3272
rect 435364 3324 435416 3330
rect 435364 3266 435416 3272
rect 433248 2984 433300 2990
rect 433248 2926 433300 2932
rect 433260 480 433288 2926
rect 434456 480 434484 3266
rect 435548 2984 435600 2990
rect 435548 2926 435600 2932
rect 435560 480 435588 2926
rect 436756 480 436784 3334
rect 437940 3324 437992 3330
rect 437940 3266 437992 3272
rect 437952 480 437980 3266
rect 439148 480 439176 3334
rect 440344 480 440372 3946
rect 440896 3330 440924 278462
rect 440884 3324 440936 3330
rect 440884 3266 440936 3272
rect 441528 3324 441580 3330
rect 441528 3266 441580 3272
rect 441540 480 441568 3266
rect 442276 2922 442304 278938
rect 442368 277914 442396 281846
rect 442356 277908 442408 277914
rect 442356 277850 442408 277856
rect 443104 3874 443132 281846
rect 443932 279070 443960 281846
rect 444288 279404 444340 279410
rect 444288 279346 444340 279352
rect 443920 279064 443972 279070
rect 443920 279006 443972 279012
rect 443092 3868 443144 3874
rect 443092 3810 443144 3816
rect 444300 3602 444328 279346
rect 444760 277982 444788 281846
rect 445772 279886 445800 281846
rect 445760 279880 445812 279886
rect 445760 279822 445812 279828
rect 446508 279002 446536 281846
rect 446496 278996 446548 279002
rect 446496 278938 446548 278944
rect 444748 277976 444800 277982
rect 444748 277918 444800 277924
rect 446404 277976 446456 277982
rect 446404 277918 446456 277924
rect 445760 6180 445812 6186
rect 445760 6122 445812 6128
rect 443828 3596 443880 3602
rect 443828 3538 443880 3544
rect 444288 3596 444340 3602
rect 444288 3538 444340 3544
rect 442632 3052 442684 3058
rect 442632 2994 442684 3000
rect 442264 2916 442316 2922
rect 442264 2858 442316 2864
rect 442644 480 442672 2994
rect 443840 480 443868 3538
rect 445772 2990 445800 6122
rect 446220 4072 446272 4078
rect 446220 4014 446272 4020
rect 445024 2984 445076 2990
rect 445024 2926 445076 2932
rect 445760 2984 445812 2990
rect 445760 2926 445812 2932
rect 445036 480 445064 2926
rect 446232 480 446260 4014
rect 446416 3330 446444 277918
rect 447336 277846 447364 281846
rect 447796 279698 447824 281846
rect 449084 280022 449112 281846
rect 449072 280016 449124 280022
rect 449072 279958 449124 279964
rect 449808 280016 449860 280022
rect 449808 279958 449860 279964
rect 447428 279670 447824 279698
rect 447324 277840 447376 277846
rect 447324 277782 447376 277788
rect 447428 277394 447456 279670
rect 449164 279200 449216 279206
rect 449164 279142 449216 279148
rect 447784 278656 447836 278662
rect 447784 278598 447836 278604
rect 447152 277366 447456 277394
rect 447152 3874 447180 277366
rect 447140 3868 447192 3874
rect 447140 3810 447192 3816
rect 446404 3324 446456 3330
rect 446404 3266 446456 3272
rect 447416 3324 447468 3330
rect 447416 3266 447468 3272
rect 447428 480 447456 3266
rect 447796 3058 447824 278598
rect 448612 3596 448664 3602
rect 448612 3538 448664 3544
rect 447784 3052 447836 3058
rect 447784 2994 447836 3000
rect 448624 480 448652 3538
rect 449176 2922 449204 279142
rect 449164 2916 449216 2922
rect 449164 2858 449216 2864
rect 449820 480 449848 279958
rect 449912 278118 449940 281846
rect 450740 279954 450768 281846
rect 450728 279948 450780 279954
rect 450728 279890 450780 279896
rect 451188 279880 451240 279886
rect 451188 279822 451240 279828
rect 449900 278112 449952 278118
rect 449900 278054 449952 278060
rect 450544 278112 450596 278118
rect 450544 278054 450596 278060
rect 450556 3602 450584 278054
rect 451200 6914 451228 279822
rect 450924 6886 451228 6914
rect 450544 3596 450596 3602
rect 450544 3538 450596 3544
rect 450924 480 450952 6886
rect 451292 4146 451320 281846
rect 452672 278050 452700 281846
rect 452660 278044 452712 278050
rect 452660 277986 452712 277992
rect 452948 277394 452976 281846
rect 454144 279614 454172 281846
rect 454684 279948 454736 279954
rect 454684 279890 454736 279896
rect 454132 279608 454184 279614
rect 454132 279550 454184 279556
rect 453304 278044 453356 278050
rect 453304 277986 453356 277992
rect 452672 277366 452976 277394
rect 451280 4140 451332 4146
rect 451280 4082 451332 4088
rect 452108 3392 452160 3398
rect 452108 3334 452160 3340
rect 452120 480 452148 3334
rect 452672 3262 452700 277366
rect 453316 3398 453344 277986
rect 453304 3392 453356 3398
rect 453304 3334 453356 3340
rect 452660 3256 452712 3262
rect 452660 3198 452712 3204
rect 453304 3256 453356 3262
rect 453304 3198 453356 3204
rect 453316 480 453344 3198
rect 454500 3052 454552 3058
rect 454500 2994 454552 3000
rect 454512 480 454540 2994
rect 454696 2854 454724 279890
rect 454776 279268 454828 279274
rect 454776 279210 454828 279216
rect 454788 3194 454816 279210
rect 455064 278186 455092 281846
rect 455892 278934 455920 281846
rect 457042 281602 457070 281860
rect 456996 281574 457070 281602
rect 457548 281846 457884 281874
rect 458468 281846 458804 281874
rect 456064 279132 456116 279138
rect 456064 279074 456116 279080
rect 455880 278928 455932 278934
rect 455880 278870 455932 278876
rect 455052 278180 455104 278186
rect 455052 278122 455104 278128
rect 456076 3466 456104 279074
rect 456892 4140 456944 4146
rect 456892 4082 456944 4088
rect 456064 3460 456116 3466
rect 456064 3402 456116 3408
rect 455696 3324 455748 3330
rect 455696 3266 455748 3272
rect 454776 3188 454828 3194
rect 454776 3130 454828 3136
rect 454684 2848 454736 2854
rect 454684 2790 454736 2796
rect 455708 480 455736 3266
rect 456904 480 456932 4082
rect 456996 3398 457024 281574
rect 457548 278254 457576 281846
rect 458088 279608 458140 279614
rect 458088 279550 458140 279556
rect 457536 278248 457588 278254
rect 457536 278190 457588 278196
rect 456984 3392 457036 3398
rect 456984 3334 457036 3340
rect 458100 480 458128 279550
rect 458468 279274 458496 281846
rect 459618 281602 459646 281860
rect 459572 281574 459646 281602
rect 460124 281846 460460 281874
rect 461044 281846 461288 281874
rect 461504 281846 462208 281874
rect 462700 281846 463036 281874
rect 463712 281846 463864 281874
rect 464356 281846 464692 281874
rect 465276 281846 465612 281874
rect 466104 281846 466440 281874
rect 466932 281846 467268 281874
rect 467852 281846 468096 281874
rect 468220 281846 469016 281874
rect 469508 281846 469844 281874
rect 459572 279478 459600 281574
rect 459560 279472 459612 279478
rect 459560 279414 459612 279420
rect 458456 279268 458508 279274
rect 458456 279210 458508 279216
rect 460124 277778 460152 281846
rect 461044 279546 461072 281846
rect 461032 279540 461084 279546
rect 461032 279482 461084 279488
rect 460296 279268 460348 279274
rect 460296 279210 460348 279216
rect 460204 279064 460256 279070
rect 460204 279006 460256 279012
rect 460112 277772 460164 277778
rect 460112 277714 460164 277720
rect 460216 4078 460244 279006
rect 460204 4072 460256 4078
rect 460204 4014 460256 4020
rect 459192 4004 459244 4010
rect 459192 3946 459244 3952
rect 459204 480 459232 3946
rect 460308 3262 460336 279210
rect 461504 277394 461532 281846
rect 461584 279336 461636 279342
rect 461584 279278 461636 279284
rect 461044 277366 461532 277394
rect 461044 3534 461072 277366
rect 461596 4146 461624 279278
rect 462700 278322 462728 281846
rect 463712 279954 463740 281846
rect 464356 280158 464384 281846
rect 464344 280152 464396 280158
rect 464344 280094 464396 280100
rect 463700 279948 463752 279954
rect 463700 279890 463752 279896
rect 464436 279540 464488 279546
rect 464436 279482 464488 279488
rect 464344 279472 464396 279478
rect 464344 279414 464396 279420
rect 462964 278928 463016 278934
rect 462964 278870 463016 278876
rect 462688 278316 462740 278322
rect 462688 278258 462740 278264
rect 461584 4140 461636 4146
rect 461584 4082 461636 4088
rect 462780 4072 462832 4078
rect 462780 4014 462832 4020
rect 461032 3528 461084 3534
rect 461032 3470 461084 3476
rect 460388 3460 460440 3466
rect 460388 3402 460440 3408
rect 460296 3256 460348 3262
rect 460296 3198 460348 3204
rect 460400 480 460428 3402
rect 461584 3392 461636 3398
rect 461584 3334 461636 3340
rect 461596 480 461624 3334
rect 462792 480 462820 4014
rect 462976 3466 463004 278870
rect 462964 3460 463016 3466
rect 462964 3402 463016 3408
rect 463976 3460 464028 3466
rect 463976 3402 464028 3408
rect 463988 480 464016 3402
rect 464356 3126 464384 279414
rect 464448 3738 464476 279482
rect 465276 278730 465304 281846
rect 466104 279546 466132 281846
rect 466368 279948 466420 279954
rect 466368 279890 466420 279896
rect 466092 279540 466144 279546
rect 466092 279482 466144 279488
rect 465264 278724 465316 278730
rect 465264 278666 465316 278672
rect 466276 278180 466328 278186
rect 466276 278122 466328 278128
rect 464436 3732 464488 3738
rect 464436 3674 464488 3680
rect 465172 3188 465224 3194
rect 465172 3130 465224 3136
rect 464344 3120 464396 3126
rect 464344 3062 464396 3068
rect 465184 480 465212 3130
rect 466288 480 466316 278122
rect 466380 3194 466408 279890
rect 466932 279478 466960 281846
rect 467104 279540 467156 279546
rect 467104 279482 467156 279488
rect 466920 279472 466972 279478
rect 466920 279414 466972 279420
rect 467116 3942 467144 279482
rect 467748 279472 467800 279478
rect 467748 279414 467800 279420
rect 467760 6914 467788 279414
rect 467852 278458 467880 281846
rect 467840 278452 467892 278458
rect 467840 278394 467892 278400
rect 468220 277394 468248 281846
rect 469508 279546 469536 281846
rect 470658 281602 470686 281860
rect 470612 281574 470686 281602
rect 471164 281846 471500 281874
rect 472084 281846 472420 281874
rect 472544 281846 473248 281874
rect 473740 281846 474076 281874
rect 474752 281846 474996 281874
rect 475488 281846 475824 281874
rect 476316 281846 476652 281874
rect 477144 281846 477480 281874
rect 478064 281846 478400 281874
rect 478892 281846 479228 281874
rect 479720 281846 480056 281874
rect 480548 281846 480884 281874
rect 481652 281846 481804 281874
rect 482296 281846 482632 281874
rect 483124 281846 483460 281874
rect 483952 281846 484288 281874
rect 484872 281846 485208 281874
rect 485792 281846 486036 281874
rect 486528 281846 486864 281874
rect 487356 281846 487692 281874
rect 469496 279540 469548 279546
rect 469496 279482 469548 279488
rect 468484 278996 468536 279002
rect 468484 278938 468536 278944
rect 467484 6886 467788 6914
rect 467852 277366 468248 277394
rect 467104 3936 467156 3942
rect 467104 3878 467156 3884
rect 466368 3188 466420 3194
rect 466368 3130 466420 3136
rect 467484 480 467512 6886
rect 467852 3670 467880 277366
rect 468496 3806 468524 278938
rect 469864 278792 469916 278798
rect 469864 278734 469916 278740
rect 468668 3936 468720 3942
rect 468668 3878 468720 3884
rect 468484 3800 468536 3806
rect 468484 3742 468536 3748
rect 467840 3664 467892 3670
rect 467840 3606 467892 3612
rect 468680 480 468708 3878
rect 469876 3874 469904 278734
rect 470612 278390 470640 281574
rect 471164 279206 471192 281846
rect 471888 280152 471940 280158
rect 471888 280094 471940 280100
rect 471152 279200 471204 279206
rect 471152 279142 471204 279148
rect 470600 278384 470652 278390
rect 470600 278326 470652 278332
rect 471244 278248 471296 278254
rect 471244 278190 471296 278196
rect 469864 3868 469916 3874
rect 469864 3810 469916 3816
rect 471060 3528 471112 3534
rect 471060 3470 471112 3476
rect 469864 3188 469916 3194
rect 469864 3130 469916 3136
rect 469876 480 469904 3130
rect 471072 480 471100 3470
rect 471256 3194 471284 278190
rect 471900 3534 471928 280094
rect 472084 280090 472112 281846
rect 472072 280084 472124 280090
rect 472072 280026 472124 280032
rect 472544 277394 472572 281846
rect 472624 280084 472676 280090
rect 472624 280026 472676 280032
rect 472084 277366 472572 277394
rect 472084 276690 472112 277366
rect 472072 276684 472124 276690
rect 472072 276626 472124 276632
rect 472636 3602 472664 280026
rect 473740 279682 473768 281846
rect 473728 279676 473780 279682
rect 473728 279618 473780 279624
rect 474752 279002 474780 281846
rect 474740 278996 474792 279002
rect 474740 278938 474792 278944
rect 475384 278928 475436 278934
rect 475384 278870 475436 278876
rect 474004 278860 474056 278866
rect 474004 278802 474056 278808
rect 472716 91792 472768 91798
rect 472716 91734 472768 91740
rect 472624 3596 472676 3602
rect 472624 3538 472676 3544
rect 471888 3528 471940 3534
rect 471888 3470 471940 3476
rect 472728 3398 472756 91734
rect 474016 4146 474044 278802
rect 474004 4140 474056 4146
rect 474004 4082 474056 4088
rect 473452 3732 473504 3738
rect 473452 3674 473504 3680
rect 472716 3392 472768 3398
rect 472716 3334 472768 3340
rect 472256 3324 472308 3330
rect 472256 3266 472308 3272
rect 471244 3188 471296 3194
rect 471244 3130 471296 3136
rect 472268 480 472296 3266
rect 473464 480 473492 3674
rect 475396 3670 475424 278870
rect 475488 278594 475516 281846
rect 476316 279138 476344 281846
rect 477144 279750 477172 281846
rect 477132 279744 477184 279750
rect 477132 279686 477184 279692
rect 476304 279132 476356 279138
rect 476304 279074 476356 279080
rect 476764 278996 476816 279002
rect 476764 278938 476816 278944
rect 475476 278588 475528 278594
rect 475476 278530 475528 278536
rect 476776 3942 476804 278938
rect 478064 278526 478092 281846
rect 478892 279818 478920 281846
rect 478880 279812 478932 279818
rect 478880 279754 478932 279760
rect 479524 279744 479576 279750
rect 479524 279686 479576 279692
rect 478144 279132 478196 279138
rect 478144 279074 478196 279080
rect 478052 278520 478104 278526
rect 478052 278462 478104 278468
rect 478156 6914 478184 279074
rect 478064 6886 478184 6914
rect 476764 3936 476816 3942
rect 476764 3878 476816 3884
rect 475384 3664 475436 3670
rect 475384 3606 475436 3612
rect 476948 3664 477000 3670
rect 476948 3606 477000 3612
rect 474556 3596 474608 3602
rect 474556 3538 474608 3544
rect 474568 480 474596 3538
rect 475752 3052 475804 3058
rect 475752 2994 475804 3000
rect 475764 480 475792 2994
rect 476960 480 476988 3606
rect 478064 3330 478092 6886
rect 479340 3936 479392 3942
rect 479340 3878 479392 3884
rect 478144 3528 478196 3534
rect 478144 3470 478196 3476
rect 478052 3324 478104 3330
rect 478052 3266 478104 3272
rect 478156 480 478184 3470
rect 479352 480 479380 3878
rect 479536 3534 479564 279686
rect 479616 279200 479668 279206
rect 479616 279142 479668 279148
rect 479524 3528 479576 3534
rect 479524 3470 479576 3476
rect 479628 3058 479656 279142
rect 479720 278798 479748 281846
rect 479708 278792 479760 278798
rect 479708 278734 479760 278740
rect 480548 277982 480576 281846
rect 480904 279676 480956 279682
rect 480904 279618 480956 279624
rect 480536 277976 480588 277982
rect 480536 277918 480588 277924
rect 480916 3942 480944 279618
rect 481652 278662 481680 281846
rect 482296 279410 482324 281846
rect 482928 279812 482980 279818
rect 482928 279754 482980 279760
rect 482284 279404 482336 279410
rect 482284 279346 482336 279352
rect 481640 278656 481692 278662
rect 481640 278598 481692 278604
rect 482284 278384 482336 278390
rect 482284 278326 482336 278332
rect 480904 3936 480956 3942
rect 480904 3878 480956 3884
rect 481732 3596 481784 3602
rect 481732 3538 481784 3544
rect 480536 3392 480588 3398
rect 480536 3334 480588 3340
rect 479616 3052 479668 3058
rect 479616 2994 479668 3000
rect 480548 480 480576 3334
rect 481744 480 481772 3538
rect 482296 3398 482324 278326
rect 482940 3602 482968 279754
rect 483124 6186 483152 281846
rect 483952 279070 483980 281846
rect 484872 280090 484900 281846
rect 484860 280084 484912 280090
rect 484860 280026 484912 280032
rect 485688 280084 485740 280090
rect 485688 280026 485740 280032
rect 483940 279064 483992 279070
rect 483940 279006 483992 279012
rect 485044 278452 485096 278458
rect 485044 278394 485096 278400
rect 484308 278316 484360 278322
rect 484308 278258 484360 278264
rect 484320 6914 484348 278258
rect 484044 6886 484348 6914
rect 483112 6180 483164 6186
rect 483112 6122 483164 6128
rect 482928 3596 482980 3602
rect 482928 3538 482980 3544
rect 482284 3392 482336 3398
rect 482284 3334 482336 3340
rect 482836 3324 482888 3330
rect 482836 3266 482888 3272
rect 482848 480 482876 3266
rect 484044 480 484072 6886
rect 485056 4010 485084 278394
rect 485044 4004 485096 4010
rect 485044 3946 485096 3952
rect 485700 3602 485728 280026
rect 485792 278118 485820 281846
rect 486528 280022 486556 281846
rect 486516 280016 486568 280022
rect 486516 279958 486568 279964
rect 487356 279886 487384 281846
rect 488598 281602 488626 281860
rect 488552 281574 488626 281602
rect 489104 281846 489440 281874
rect 490024 281846 490268 281874
rect 490576 281846 491096 281874
rect 491680 281846 492016 281874
rect 492692 281846 492844 281874
rect 493520 281846 493672 281874
rect 494164 281846 494500 281874
rect 495084 281846 495420 281874
rect 495912 281846 496248 281874
rect 487344 279880 487396 279886
rect 487344 279822 487396 279828
rect 487068 279404 487120 279410
rect 487068 279346 487120 279352
rect 486424 278520 486476 278526
rect 486424 278462 486476 278468
rect 485780 278112 485832 278118
rect 485780 278054 485832 278060
rect 486436 6914 486464 278462
rect 486344 6886 486464 6914
rect 486344 4078 486372 6886
rect 486332 4072 486384 4078
rect 486332 4014 486384 4020
rect 487080 3602 487108 279346
rect 488552 278050 488580 281574
rect 489104 279274 489132 281846
rect 489828 279880 489880 279886
rect 489828 279822 489880 279828
rect 489092 279268 489144 279274
rect 489092 279210 489144 279216
rect 489184 278112 489236 278118
rect 489184 278054 489236 278060
rect 488540 278044 488592 278050
rect 488540 277986 488592 277992
rect 489196 3602 489224 278054
rect 485228 3596 485280 3602
rect 485228 3538 485280 3544
rect 485688 3596 485740 3602
rect 485688 3538 485740 3544
rect 486424 3596 486476 3602
rect 486424 3538 486476 3544
rect 487068 3596 487120 3602
rect 487068 3538 487120 3544
rect 487620 3596 487672 3602
rect 487620 3538 487672 3544
rect 489184 3596 489236 3602
rect 489184 3538 489236 3544
rect 485240 480 485268 3538
rect 486436 480 486464 3538
rect 487632 480 487660 3538
rect 489840 3398 489868 279822
rect 490024 278866 490052 281846
rect 490012 278860 490064 278866
rect 490012 278802 490064 278808
rect 490576 277394 490604 281846
rect 491680 279342 491708 281846
rect 492692 279614 492720 281846
rect 492680 279608 492732 279614
rect 492680 279550 492732 279556
rect 493324 279608 493376 279614
rect 493324 279550 493376 279556
rect 491668 279336 491720 279342
rect 491668 279278 491720 279284
rect 491208 278044 491260 278050
rect 491208 277986 491260 277992
rect 490024 277366 490604 277394
rect 490024 91798 490052 277366
rect 490012 91792 490064 91798
rect 490012 91734 490064 91740
rect 491220 6914 491248 277986
rect 491128 6886 491248 6914
rect 488816 3392 488868 3398
rect 488816 3334 488868 3340
rect 489828 3392 489880 3398
rect 489828 3334 489880 3340
rect 488828 480 488856 3334
rect 489920 2984 489972 2990
rect 489920 2926 489972 2932
rect 489932 480 489960 2926
rect 491128 480 491156 6886
rect 493336 3466 493364 279550
rect 493520 278526 493548 281846
rect 494164 279546 494192 281846
rect 494152 279540 494204 279546
rect 494152 279482 494204 279488
rect 495084 278934 495112 281846
rect 495348 279540 495400 279546
rect 495348 279482 495400 279488
rect 495072 278928 495124 278934
rect 495072 278870 495124 278876
rect 493508 278520 493560 278526
rect 493508 278462 493560 278468
rect 493416 278452 493468 278458
rect 493416 278394 493468 278400
rect 493428 3738 493456 278394
rect 493508 3800 493560 3806
rect 493508 3742 493560 3748
rect 493416 3732 493468 3738
rect 493416 3674 493468 3680
rect 492312 3460 492364 3466
rect 492312 3402 492364 3408
rect 493324 3460 493376 3466
rect 493324 3402 493376 3408
rect 492324 480 492352 3402
rect 493520 480 493548 3742
rect 495360 3466 495388 279482
rect 495912 278594 495940 281846
rect 497062 281602 497090 281860
rect 497016 281574 497090 281602
rect 497660 281846 497996 281874
rect 498488 281846 498824 281874
rect 496728 280016 496780 280022
rect 496728 279958 496780 279964
rect 495900 278588 495952 278594
rect 495900 278530 495952 278536
rect 496740 3466 496768 279958
rect 494704 3460 494756 3466
rect 494704 3402 494756 3408
rect 495348 3460 495400 3466
rect 495348 3402 495400 3408
rect 495900 3460 495952 3466
rect 495900 3402 495952 3408
rect 496728 3460 496780 3466
rect 496728 3402 496780 3408
rect 494716 480 494744 3402
rect 495912 480 495940 3402
rect 497016 3398 497044 281574
rect 497660 279954 497688 281846
rect 497648 279948 497700 279954
rect 497648 279890 497700 279896
rect 497464 279064 497516 279070
rect 497464 279006 497516 279012
rect 497096 4140 497148 4146
rect 497096 4082 497148 4088
rect 497004 3392 497056 3398
rect 497004 3334 497056 3340
rect 497108 480 497136 4082
rect 497476 2990 497504 279006
rect 498488 278186 498516 281846
rect 499638 281602 499666 281860
rect 499592 281574 499666 281602
rect 500144 281846 500480 281874
rect 501064 281846 501400 281874
rect 501892 281846 502228 281874
rect 502720 281846 503056 281874
rect 503732 281846 503884 281874
rect 504008 281846 504804 281874
rect 505296 281846 505632 281874
rect 506124 281846 506460 281874
rect 506952 281846 507288 281874
rect 507872 281846 508208 281874
rect 508700 281846 509036 281874
rect 509528 281846 509864 281874
rect 499592 279478 499620 281574
rect 499580 279472 499632 279478
rect 499580 279414 499632 279420
rect 500144 279002 500172 281846
rect 500868 279472 500920 279478
rect 500868 279414 500920 279420
rect 500132 278996 500184 279002
rect 500132 278938 500184 278944
rect 498476 278180 498528 278186
rect 498476 278122 498528 278128
rect 500880 6914 500908 279414
rect 501064 278254 501092 281846
rect 501892 280158 501920 281846
rect 501880 280152 501932 280158
rect 501880 280094 501932 280100
rect 502248 279948 502300 279954
rect 502248 279890 502300 279896
rect 501604 279336 501656 279342
rect 501604 279278 501656 279284
rect 501052 278248 501104 278254
rect 501052 278190 501104 278196
rect 500604 6886 500908 6914
rect 498200 3732 498252 3738
rect 498200 3674 498252 3680
rect 497464 2984 497516 2990
rect 497464 2926 497516 2932
rect 498212 480 498240 3674
rect 499396 3460 499448 3466
rect 499396 3402 499448 3408
rect 499408 480 499436 3402
rect 500604 480 500632 6886
rect 501616 4146 501644 279278
rect 501604 4140 501656 4146
rect 501604 4082 501656 4088
rect 502260 3534 502288 279890
rect 502720 279138 502748 281846
rect 503628 280152 503680 280158
rect 503628 280094 503680 280100
rect 502984 279268 503036 279274
rect 502984 279210 503036 279216
rect 502708 279132 502760 279138
rect 502708 279074 502760 279080
rect 502996 6914 503024 279210
rect 502904 6886 503024 6914
rect 502904 3670 502932 6886
rect 502892 3664 502944 3670
rect 502892 3606 502944 3612
rect 503640 3534 503668 280094
rect 503732 278458 503760 281846
rect 503720 278452 503772 278458
rect 503720 278394 503772 278400
rect 504008 277394 504036 281846
rect 505296 279206 505324 281846
rect 506124 279274 506152 281846
rect 506952 279750 506980 281846
rect 506940 279744 506992 279750
rect 506940 279686 506992 279692
rect 507768 279744 507820 279750
rect 507768 279686 507820 279692
rect 506112 279268 506164 279274
rect 506112 279210 506164 279216
rect 505284 279200 505336 279206
rect 505284 279142 505336 279148
rect 504364 279132 504416 279138
rect 504364 279074 504416 279080
rect 503732 277366 504036 277394
rect 503732 3738 503760 277366
rect 504180 3868 504232 3874
rect 504180 3810 504232 3816
rect 503720 3732 503772 3738
rect 503720 3674 503772 3680
rect 501788 3528 501840 3534
rect 501788 3470 501840 3476
rect 502248 3528 502300 3534
rect 502248 3470 502300 3476
rect 502984 3528 503036 3534
rect 502984 3470 503036 3476
rect 503628 3528 503680 3534
rect 503628 3470 503680 3476
rect 501800 480 501828 3470
rect 502996 480 503024 3470
rect 504192 480 504220 3810
rect 504376 3806 504404 279074
rect 504364 3800 504416 3806
rect 504364 3742 504416 3748
rect 505376 3596 505428 3602
rect 505376 3538 505428 3544
rect 505388 480 505416 3538
rect 507676 3528 507728 3534
rect 507676 3470 507728 3476
rect 506480 3256 506532 3262
rect 506480 3198 506532 3204
rect 506492 480 506520 3198
rect 507688 480 507716 3470
rect 507780 3262 507808 279686
rect 507872 279682 507900 281846
rect 507860 279676 507912 279682
rect 507860 279618 507912 279624
rect 508504 278996 508556 279002
rect 508504 278938 508556 278944
rect 508516 3942 508544 278938
rect 508700 278390 508728 281846
rect 509528 279818 509556 281846
rect 510678 281602 510706 281860
rect 510632 281574 510706 281602
rect 511276 281846 511612 281874
rect 512104 281846 512440 281874
rect 512932 281846 513268 281874
rect 513760 281846 514096 281874
rect 514772 281846 515016 281874
rect 515508 281846 515844 281874
rect 516336 281846 516672 281874
rect 509516 279812 509568 279818
rect 509516 279754 509568 279760
rect 509148 279676 509200 279682
rect 509148 279618 509200 279624
rect 508688 278384 508740 278390
rect 508688 278326 508740 278332
rect 509160 6914 509188 279618
rect 508884 6886 509188 6914
rect 508504 3936 508556 3942
rect 508504 3878 508556 3884
rect 507768 3256 507820 3262
rect 507768 3198 507820 3204
rect 508884 480 508912 6886
rect 510632 3670 510660 281574
rect 511276 278322 511304 281846
rect 512104 280090 512132 281846
rect 512092 280084 512144 280090
rect 512092 280026 512144 280032
rect 512932 279410 512960 281846
rect 513288 280084 513340 280090
rect 513288 280026 513340 280032
rect 512920 279404 512972 279410
rect 512920 279346 512972 279352
rect 511908 279268 511960 279274
rect 511908 279210 511960 279216
rect 511264 278316 511316 278322
rect 511264 278258 511316 278264
rect 510620 3664 510672 3670
rect 510620 3606 510672 3612
rect 511920 3466 511948 279210
rect 512644 278928 512696 278934
rect 512644 278870 512696 278876
rect 512656 3874 512684 278870
rect 512644 3868 512696 3874
rect 512644 3810 512696 3816
rect 513300 3466 513328 280026
rect 513760 278118 513788 281846
rect 514772 279886 514800 281846
rect 514760 279880 514812 279886
rect 514760 279822 514812 279828
rect 514668 279812 514720 279818
rect 514668 279754 514720 279760
rect 513748 278112 513800 278118
rect 513748 278054 513800 278060
rect 514680 3466 514708 279754
rect 515508 279070 515536 281846
rect 516048 279880 516100 279886
rect 516048 279822 516100 279828
rect 515956 279404 516008 279410
rect 515956 279346 516008 279352
rect 515496 279064 515548 279070
rect 515496 279006 515548 279012
rect 515968 16574 515996 279346
rect 515876 16546 515996 16574
rect 515876 3466 515904 16546
rect 516060 6914 516088 279822
rect 516336 278050 516364 281846
rect 517578 281602 517606 281860
rect 517532 281574 517606 281602
rect 518084 281846 518420 281874
rect 518912 281846 519248 281874
rect 519740 281846 520076 281874
rect 520660 281846 520996 281874
rect 521672 281846 521824 281874
rect 521948 281846 522652 281874
rect 523144 281846 523480 281874
rect 524064 281846 524400 281874
rect 524892 281846 525228 281874
rect 525812 281846 526056 281874
rect 526548 281846 526884 281874
rect 527468 281846 527804 281874
rect 517532 279614 517560 281574
rect 517520 279608 517572 279614
rect 517520 279550 517572 279556
rect 517428 279200 517480 279206
rect 517428 279142 517480 279148
rect 516324 278044 516376 278050
rect 516324 277986 516376 277992
rect 517440 6914 517468 279142
rect 518084 279138 518112 281846
rect 518912 279546 518940 281846
rect 519740 280022 519768 281846
rect 519728 280016 519780 280022
rect 519728 279958 519780 279964
rect 519544 279744 519596 279750
rect 519544 279686 519596 279692
rect 518900 279540 518952 279546
rect 518900 279482 518952 279488
rect 518072 279132 518124 279138
rect 518072 279074 518124 279080
rect 518164 279132 518216 279138
rect 518164 279074 518216 279080
rect 515968 6886 516088 6914
rect 517164 6886 517468 6914
rect 511264 3460 511316 3466
rect 511264 3402 511316 3408
rect 511908 3460 511960 3466
rect 511908 3402 511960 3408
rect 512460 3460 512512 3466
rect 512460 3402 512512 3408
rect 513288 3460 513340 3466
rect 513288 3402 513340 3408
rect 513564 3460 513616 3466
rect 513564 3402 513616 3408
rect 514668 3460 514720 3466
rect 514668 3402 514720 3408
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 515864 3460 515916 3466
rect 515864 3402 515916 3408
rect 510068 3324 510120 3330
rect 510068 3266 510120 3272
rect 510080 480 510108 3266
rect 511276 480 511304 3402
rect 512472 480 512500 3402
rect 513576 480 513604 3402
rect 514772 480 514800 3402
rect 515968 480 515996 6886
rect 517164 480 517192 6886
rect 518176 3330 518204 279074
rect 519556 3670 519584 279686
rect 520188 279540 520240 279546
rect 520188 279482 520240 279488
rect 519544 3664 519596 3670
rect 519544 3606 519596 3612
rect 518348 3596 518400 3602
rect 518348 3538 518400 3544
rect 518164 3324 518216 3330
rect 518164 3266 518216 3272
rect 518360 480 518388 3538
rect 520200 3466 520228 279482
rect 520660 279342 520688 281846
rect 520648 279336 520700 279342
rect 520648 279278 520700 279284
rect 521568 279064 521620 279070
rect 521568 279006 521620 279012
rect 521580 3466 521608 279006
rect 521672 279002 521700 281846
rect 521660 278996 521712 279002
rect 521660 278938 521712 278944
rect 519544 3460 519596 3466
rect 519544 3402 519596 3408
rect 520188 3460 520240 3466
rect 520188 3402 520240 3408
rect 520740 3460 520792 3466
rect 520740 3402 520792 3408
rect 521568 3460 521620 3466
rect 521568 3402 521620 3408
rect 521844 3460 521896 3466
rect 521844 3402 521896 3408
rect 519556 480 519584 3402
rect 520752 480 520780 3402
rect 521856 480 521884 3402
rect 521948 3398 521976 281846
rect 522948 279608 523000 279614
rect 522948 279550 523000 279556
rect 522960 3466 522988 279550
rect 523144 279478 523172 281846
rect 524064 279954 524092 281846
rect 524892 280158 524920 281846
rect 524880 280152 524932 280158
rect 524880 280094 524932 280100
rect 525156 280152 525208 280158
rect 525156 280094 525208 280100
rect 524052 279948 524104 279954
rect 524052 279890 524104 279896
rect 525064 279948 525116 279954
rect 525064 279890 525116 279896
rect 523132 279472 523184 279478
rect 523132 279414 523184 279420
rect 522948 3460 523000 3466
rect 522948 3402 523000 3408
rect 524236 3460 524288 3466
rect 524236 3402 524288 3408
rect 521936 3392 521988 3398
rect 521936 3334 521988 3340
rect 523040 3392 523092 3398
rect 523040 3334 523092 3340
rect 523052 480 523080 3334
rect 524248 480 524276 3402
rect 525076 3398 525104 279890
rect 525168 3466 525196 280094
rect 525812 278934 525840 281846
rect 526548 279750 526576 281846
rect 527468 280022 527496 281846
rect 528618 281602 528646 281860
rect 529124 281846 529460 281874
rect 529952 281846 530288 281874
rect 530872 281846 531208 281874
rect 531700 281846 532036 281874
rect 532712 281846 532864 281874
rect 533540 281846 533692 281874
rect 534276 281846 534612 281874
rect 535104 281846 535440 281874
rect 535564 281846 536268 281874
rect 536852 281846 537096 281874
rect 537680 281846 538016 281874
rect 538508 281846 538844 281874
rect 528618 281574 528692 281602
rect 527456 280016 527508 280022
rect 527456 279958 527508 279964
rect 526536 279744 526588 279750
rect 526536 279686 526588 279692
rect 526444 279472 526496 279478
rect 526444 279414 526496 279420
rect 525800 278928 525852 278934
rect 525800 278870 525852 278876
rect 525156 3460 525208 3466
rect 525156 3402 525208 3408
rect 525064 3392 525116 3398
rect 525064 3334 525116 3340
rect 526456 2990 526484 279414
rect 527088 279336 527140 279342
rect 527088 279278 527140 279284
rect 527100 3466 527128 279278
rect 528664 3534 528692 281574
rect 529124 279682 529152 281846
rect 529112 279676 529164 279682
rect 529112 279618 529164 279624
rect 529848 279676 529900 279682
rect 529848 279618 529900 279624
rect 529860 3534 529888 279618
rect 529952 279138 529980 281846
rect 530872 279274 530900 281846
rect 531700 280090 531728 281846
rect 531688 280084 531740 280090
rect 531688 280026 531740 280032
rect 532712 279818 532740 281846
rect 533436 280084 533488 280090
rect 533436 280026 533488 280032
rect 532700 279812 532752 279818
rect 532700 279754 532752 279760
rect 533344 279812 533396 279818
rect 533344 279754 533396 279760
rect 530860 279268 530912 279274
rect 530860 279210 530912 279216
rect 531228 279268 531280 279274
rect 531228 279210 531280 279216
rect 529940 279132 529992 279138
rect 529940 279074 529992 279080
rect 528652 3528 528704 3534
rect 528652 3470 528704 3476
rect 529020 3528 529072 3534
rect 529020 3470 529072 3476
rect 529848 3528 529900 3534
rect 529848 3470 529900 3476
rect 526628 3460 526680 3466
rect 526628 3402 526680 3408
rect 527088 3460 527140 3466
rect 527088 3402 527140 3408
rect 527824 3460 527876 3466
rect 527824 3402 527876 3408
rect 525432 2984 525484 2990
rect 525432 2926 525484 2932
rect 526444 2984 526496 2990
rect 526444 2926 526496 2932
rect 525444 480 525472 2926
rect 526640 480 526668 3402
rect 527836 480 527864 3402
rect 529032 480 529060 3470
rect 531240 3194 531268 279210
rect 533356 3534 533384 279754
rect 532516 3528 532568 3534
rect 532516 3470 532568 3476
rect 533344 3528 533396 3534
rect 533344 3470 533396 3476
rect 531320 3392 531372 3398
rect 531320 3334 531372 3340
rect 530124 3188 530176 3194
rect 530124 3130 530176 3136
rect 531228 3188 531280 3194
rect 531228 3130 531280 3136
rect 530136 480 530164 3130
rect 531332 480 531360 3334
rect 532528 480 532556 3470
rect 533448 3398 533476 280026
rect 533540 279410 533568 281846
rect 534276 279886 534304 281846
rect 534264 279880 534316 279886
rect 534264 279822 534316 279828
rect 533528 279404 533580 279410
rect 533528 279346 533580 279352
rect 535104 279206 535132 281846
rect 535368 279744 535420 279750
rect 535368 279686 535420 279692
rect 535092 279200 535144 279206
rect 535092 279142 535144 279148
rect 533712 3596 533764 3602
rect 533712 3538 533764 3544
rect 533436 3392 533488 3398
rect 533436 3334 533488 3340
rect 533724 480 533752 3538
rect 535380 3534 535408 279686
rect 535564 3670 535592 281846
rect 536748 279880 536800 279886
rect 536748 279822 536800 279828
rect 535552 3664 535604 3670
rect 535552 3606 535604 3612
rect 536760 3534 536788 279822
rect 536852 279546 536880 281846
rect 537680 280022 537708 281846
rect 537668 280016 537720 280022
rect 537668 279958 537720 279964
rect 538128 280016 538180 280022
rect 538128 279958 538180 279964
rect 536840 279540 536892 279546
rect 536840 279482 536892 279488
rect 538140 3534 538168 279958
rect 538508 279614 538536 281846
rect 539658 281602 539686 281860
rect 539612 281574 539686 281602
rect 540256 281846 540592 281874
rect 541084 281846 541420 281874
rect 541912 281846 542248 281874
rect 542372 281846 543076 281874
rect 543752 281846 543996 281874
rect 544488 281846 544824 281874
rect 545316 281846 545652 281874
rect 546144 281846 546480 281874
rect 546696 281846 547400 281874
rect 548076 281846 548228 281874
rect 548720 281846 549056 281874
rect 549548 281846 549884 281874
rect 550652 281846 550804 281874
rect 550928 281846 551632 281874
rect 552124 281846 552460 281874
rect 552952 281846 553288 281874
rect 553872 281846 554208 281874
rect 554792 281846 555036 281874
rect 555528 281846 555864 281874
rect 556356 281846 556692 281874
rect 539612 279954 539640 281574
rect 540256 280158 540284 281846
rect 540244 280152 540296 280158
rect 540244 280094 540296 280100
rect 539600 279948 539652 279954
rect 539600 279890 539652 279896
rect 538496 279608 538548 279614
rect 538496 279550 538548 279556
rect 539508 279608 539560 279614
rect 539508 279550 539560 279556
rect 539520 3534 539548 279550
rect 540888 279540 540940 279546
rect 540888 279482 540940 279488
rect 540900 6914 540928 279482
rect 541084 279478 541112 281846
rect 541072 279472 541124 279478
rect 541072 279414 541124 279420
rect 541912 279342 541940 281846
rect 541900 279336 541952 279342
rect 541900 279278 541952 279284
rect 540808 6886 540928 6914
rect 539600 3732 539652 3738
rect 539600 3674 539652 3680
rect 534908 3528 534960 3534
rect 534908 3470 534960 3476
rect 535368 3528 535420 3534
rect 535368 3470 535420 3476
rect 536104 3528 536156 3534
rect 536104 3470 536156 3476
rect 536748 3528 536800 3534
rect 536748 3470 536800 3476
rect 537208 3528 537260 3534
rect 537208 3470 537260 3476
rect 538128 3528 538180 3534
rect 538128 3470 538180 3476
rect 538404 3528 538456 3534
rect 538404 3470 538456 3476
rect 539508 3528 539560 3534
rect 539508 3470 539560 3476
rect 534920 480 534948 3470
rect 536116 480 536144 3470
rect 537220 480 537248 3470
rect 538416 480 538444 3470
rect 539612 480 539640 3674
rect 540808 480 540836 6886
rect 541992 3528 542044 3534
rect 541992 3470 542044 3476
rect 542004 480 542032 3470
rect 542372 3466 542400 281846
rect 543004 279948 543056 279954
rect 543004 279890 543056 279896
rect 543016 3534 543044 279890
rect 543752 279682 543780 281846
rect 543740 279676 543792 279682
rect 543740 279618 543792 279624
rect 544384 279676 544436 279682
rect 544384 279618 544436 279624
rect 544396 6914 544424 279618
rect 544488 279274 544516 281846
rect 545316 280090 545344 281846
rect 545304 280084 545356 280090
rect 545304 280026 545356 280032
rect 546144 279818 546172 281846
rect 546132 279812 546184 279818
rect 546132 279754 546184 279760
rect 545028 279472 545080 279478
rect 545028 279414 545080 279420
rect 544476 279268 544528 279274
rect 544476 279210 544528 279216
rect 544304 6886 544424 6914
rect 544304 3534 544332 6886
rect 545040 3534 545068 279414
rect 546696 6914 546724 281846
rect 547144 279812 547196 279818
rect 547144 279754 547196 279760
rect 546604 6886 546724 6914
rect 546604 3602 546632 6886
rect 546592 3596 546644 3602
rect 546592 3538 546644 3544
rect 546684 3596 546736 3602
rect 546684 3538 546736 3544
rect 543004 3528 543056 3534
rect 543004 3470 543056 3476
rect 543188 3528 543240 3534
rect 543188 3470 543240 3476
rect 544292 3528 544344 3534
rect 544292 3470 544344 3476
rect 544384 3528 544436 3534
rect 544384 3470 544436 3476
rect 545028 3528 545080 3534
rect 545028 3470 545080 3476
rect 545488 3528 545540 3534
rect 545488 3470 545540 3476
rect 542360 3460 542412 3466
rect 542360 3402 542412 3408
rect 543200 480 543228 3470
rect 544396 480 544424 3470
rect 545500 480 545528 3470
rect 546696 480 546724 3538
rect 547156 3534 547184 279754
rect 548076 279750 548104 281846
rect 548720 279886 548748 281846
rect 549548 280022 549576 281846
rect 549536 280016 549588 280022
rect 549536 279958 549588 279964
rect 548708 279880 548760 279886
rect 548708 279822 548760 279828
rect 548064 279744 548116 279750
rect 548064 279686 548116 279692
rect 549168 279744 549220 279750
rect 549168 279686 549220 279692
rect 548524 279268 548576 279274
rect 548524 279210 548576 279216
rect 548536 3602 548564 279210
rect 549180 6914 549208 279686
rect 550652 279614 550680 281846
rect 550640 279608 550692 279614
rect 550640 279550 550692 279556
rect 549088 6886 549208 6914
rect 548524 3596 548576 3602
rect 548524 3538 548576 3544
rect 547144 3528 547196 3534
rect 547144 3470 547196 3476
rect 547880 3052 547932 3058
rect 547880 2994 547932 3000
rect 547892 480 547920 2994
rect 549088 480 549116 6886
rect 550928 3738 550956 281846
rect 552124 279546 552152 281846
rect 552952 279954 552980 281846
rect 552940 279948 552992 279954
rect 552940 279890 552992 279896
rect 553872 279682 553900 281846
rect 553860 279676 553912 279682
rect 553860 279618 553912 279624
rect 552112 279540 552164 279546
rect 552112 279482 552164 279488
rect 554688 279540 554740 279546
rect 554688 279482 554740 279488
rect 551284 278928 551336 278934
rect 551284 278870 551336 278876
rect 550916 3732 550968 3738
rect 550916 3674 550968 3680
rect 551296 3534 551324 278870
rect 551468 3596 551520 3602
rect 551468 3538 551520 3544
rect 550272 3528 550324 3534
rect 550272 3470 550324 3476
rect 551284 3528 551336 3534
rect 551284 3470 551336 3476
rect 550284 480 550312 3470
rect 551480 480 551508 3538
rect 554700 3534 554728 279482
rect 554792 279478 554820 281846
rect 555528 279818 555556 281846
rect 555516 279812 555568 279818
rect 555516 279754 555568 279760
rect 554780 279472 554832 279478
rect 554780 279414 554832 279420
rect 556356 279274 556384 281846
rect 557598 281602 557626 281860
rect 557552 281574 557626 281602
rect 558104 281846 558440 281874
rect 558932 281846 559268 281874
rect 559760 281846 560096 281874
rect 560404 281846 561016 281874
rect 561692 281846 561844 281874
rect 562336 281846 562672 281874
rect 563256 281846 563592 281874
rect 564084 281846 564420 281874
rect 564636 281846 565248 281874
rect 557448 279472 557500 279478
rect 557448 279414 557500 279420
rect 556344 279268 556396 279274
rect 556344 279210 556396 279216
rect 556804 278860 556856 278866
rect 556804 278802 556856 278808
rect 555424 278792 555476 278798
rect 555424 278734 555476 278740
rect 554964 3664 555016 3670
rect 554964 3606 555016 3612
rect 553768 3528 553820 3534
rect 553768 3470 553820 3476
rect 554688 3528 554740 3534
rect 554688 3470 554740 3476
rect 552664 3460 552716 3466
rect 552664 3402 552716 3408
rect 552676 480 552704 3402
rect 553780 480 553808 3470
rect 554976 480 555004 3606
rect 555436 3058 555464 278734
rect 556160 4140 556212 4146
rect 556160 4082 556212 4088
rect 555424 3052 555476 3058
rect 555424 2994 555476 3000
rect 556172 480 556200 4082
rect 556816 3602 556844 278802
rect 557460 6914 557488 279414
rect 557552 278798 557580 281574
rect 558104 279750 558132 281846
rect 558092 279744 558144 279750
rect 558092 279686 558144 279692
rect 558184 279676 558236 279682
rect 558184 279618 558236 279624
rect 557540 278792 557592 278798
rect 557540 278734 557592 278740
rect 557368 6886 557488 6914
rect 556804 3596 556856 3602
rect 556804 3538 556856 3544
rect 557368 480 557396 6886
rect 558196 3670 558224 279618
rect 558276 279608 558328 279614
rect 558276 279550 558328 279556
rect 558288 4146 558316 279550
rect 558932 278934 558960 281846
rect 558920 278928 558972 278934
rect 558920 278870 558972 278876
rect 559760 278866 559788 281846
rect 559748 278860 559800 278866
rect 559748 278802 559800 278808
rect 558276 4140 558328 4146
rect 558276 4082 558328 4088
rect 558184 3664 558236 3670
rect 558184 3606 558236 3612
rect 559748 3596 559800 3602
rect 559748 3538 559800 3544
rect 558552 3052 558604 3058
rect 558552 2994 558604 3000
rect 558564 480 558592 2994
rect 559760 480 559788 3538
rect 560404 3466 560432 281846
rect 561692 279546 561720 281846
rect 562336 279682 562364 281846
rect 562324 279676 562376 279682
rect 562324 279618 562376 279624
rect 563256 279614 563284 281846
rect 563244 279608 563296 279614
rect 563244 279550 563296 279556
rect 561680 279540 561732 279546
rect 561680 279482 561732 279488
rect 564084 279478 564112 281846
rect 564072 279472 564124 279478
rect 564072 279414 564124 279420
rect 561588 279268 561640 279274
rect 561588 279210 561640 279216
rect 561600 3534 561628 279210
rect 562968 278860 563020 278866
rect 562968 278802 563020 278808
rect 562980 3534 563008 278802
rect 563244 4004 563296 4010
rect 563244 3946 563296 3952
rect 560852 3528 560904 3534
rect 560852 3470 560904 3476
rect 561588 3528 561640 3534
rect 561588 3470 561640 3476
rect 562048 3528 562100 3534
rect 562048 3470 562100 3476
rect 562968 3528 563020 3534
rect 562968 3470 563020 3476
rect 560392 3460 560444 3466
rect 560392 3402 560444 3408
rect 560864 480 560892 3470
rect 562060 480 562088 3470
rect 563256 480 563284 3946
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564452 480 564480 3470
rect 564636 3058 564664 281846
rect 566062 281602 566090 281860
rect 566016 281574 566090 281602
rect 566660 281846 566996 281874
rect 567488 281846 567824 281874
rect 565728 279472 565780 279478
rect 565728 279414 565780 279420
rect 565740 6914 565768 279414
rect 565648 6886 565768 6914
rect 564624 3052 564676 3058
rect 564624 2994 564676 3000
rect 565648 480 565676 6886
rect 566016 3602 566044 281574
rect 566660 279274 566688 281846
rect 566648 279268 566700 279274
rect 566648 279210 566700 279216
rect 567488 278866 567516 281846
rect 568638 281602 568666 281860
rect 568592 281574 568666 281602
rect 569144 281846 569480 281874
rect 570064 281846 570400 281874
rect 570616 281846 571228 281874
rect 571720 281846 572056 281874
rect 567476 278860 567528 278866
rect 567476 278802 567528 278808
rect 566464 278792 566516 278798
rect 566464 278734 566516 278740
rect 566004 3596 566056 3602
rect 566004 3538 566056 3544
rect 566476 3534 566504 278734
rect 568592 4010 568620 281574
rect 569144 278798 569172 281846
rect 569224 279540 569276 279546
rect 569224 279482 569276 279488
rect 569132 278792 569184 278798
rect 569132 278734 569184 278740
rect 568580 4004 568632 4010
rect 568580 3946 568632 3952
rect 566832 3664 566884 3670
rect 566832 3606 566884 3612
rect 566464 3528 566516 3534
rect 566464 3470 566516 3476
rect 566844 480 566872 3606
rect 569236 3534 569264 279482
rect 570064 279478 570092 281846
rect 570052 279472 570104 279478
rect 570052 279414 570104 279420
rect 570616 277394 570644 281846
rect 571720 279546 571748 281846
rect 572870 281602 572898 281860
rect 572824 281574 572898 281602
rect 573468 281846 573804 281874
rect 574296 281846 574632 281874
rect 574848 281846 575460 281874
rect 575584 281846 576288 281874
rect 576964 281846 577208 281874
rect 577700 281846 578036 281874
rect 578252 281846 578864 281874
rect 572720 279676 572772 279682
rect 572720 279618 572772 279624
rect 572628 279608 572680 279614
rect 572628 279550 572680 279556
rect 571708 279540 571760 279546
rect 571708 279482 571760 279488
rect 570156 277366 570644 277394
rect 570156 3670 570184 277366
rect 570144 3664 570196 3670
rect 570144 3606 570196 3612
rect 570328 3596 570380 3602
rect 570328 3538 570380 3544
rect 568028 3528 568080 3534
rect 568028 3470 568080 3476
rect 569224 3528 569276 3534
rect 569224 3470 569276 3476
rect 568040 480 568068 3470
rect 569132 3188 569184 3194
rect 569132 3130 569184 3136
rect 569144 480 569172 3130
rect 570340 480 570368 3538
rect 572640 3534 572668 279550
rect 572732 3602 572760 279618
rect 572824 16574 572852 281574
rect 573468 279682 573496 281846
rect 573456 279676 573508 279682
rect 573456 279618 573508 279624
rect 574296 279614 574324 281846
rect 574284 279608 574336 279614
rect 574284 279550 574336 279556
rect 574848 277394 574876 281846
rect 575388 278792 575440 278798
rect 575388 278734 575440 278740
rect 574204 277366 574876 277394
rect 572824 16546 572944 16574
rect 572720 3596 572772 3602
rect 572720 3538 572772 3544
rect 571524 3528 571576 3534
rect 571524 3470 571576 3476
rect 572628 3528 572680 3534
rect 572628 3470 572680 3476
rect 571536 480 571564 3470
rect 572916 3194 572944 16546
rect 572904 3188 572956 3194
rect 572904 3130 572956 3136
rect 573916 3120 573968 3126
rect 573916 3062 573968 3068
rect 572720 2984 572772 2990
rect 572720 2926 572772 2932
rect 572732 480 572760 2926
rect 573928 480 573956 3062
rect 574204 2990 574232 277366
rect 575400 6914 575428 278734
rect 575124 6886 575428 6914
rect 574192 2984 574244 2990
rect 574192 2926 574244 2932
rect 575124 480 575152 6886
rect 575584 3126 575612 281846
rect 576860 280154 576912 280158
rect 576780 280152 576912 280154
rect 576780 280126 576860 280152
rect 576780 3466 576808 280126
rect 576860 280094 576912 280100
rect 576964 278798 576992 281846
rect 577700 280158 577728 281846
rect 577688 280152 577740 280158
rect 577688 280094 577740 280100
rect 576952 278792 577004 278798
rect 576952 278734 577004 278740
rect 578252 3534 578280 281846
rect 579678 281602 579706 281860
rect 579632 281574 579706 281602
rect 577412 3528 577464 3534
rect 577412 3470 577464 3476
rect 578240 3528 578292 3534
rect 578240 3470 578292 3476
rect 576308 3460 576360 3466
rect 576308 3402 576360 3408
rect 576768 3460 576820 3466
rect 576768 3402 576820 3408
rect 575572 3120 575624 3126
rect 575572 3062 575624 3068
rect 576320 480 576348 3402
rect 577424 480 577452 3470
rect 579632 3058 579660 281574
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 579988 219428 580040 219434
rect 579988 219370 580040 219376
rect 580000 219065 580028 219370
rect 579986 219056 580042 219065
rect 579986 218991 580042 219000
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 579896 60716 579948 60722
rect 579896 60658 579948 60664
rect 579908 59673 579936 60658
rect 579894 59664 579950 59673
rect 579894 59599 579950 59608
rect 580276 46345 580304 282270
rect 580356 282260 580408 282266
rect 580356 282202 580408 282208
rect 580368 73001 580396 282202
rect 580448 282192 580500 282198
rect 580448 282134 580500 282140
rect 580460 86193 580488 282134
rect 580612 281846 580856 281874
rect 580446 86184 580502 86193
rect 580446 86119 580502 86128
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580262 46336 580318 46345
rect 580262 46271 580318 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 580828 16574 580856 281846
rect 581196 281846 581440 281874
rect 581196 16574 581224 281846
rect 582254 281602 582282 281860
rect 582254 281574 582328 281602
rect 582300 279682 582328 281574
rect 582288 279676 582340 279682
rect 582288 279618 582340 279624
rect 582392 139369 582420 700159
rect 582484 152697 582512 701655
rect 582576 232393 582604 701791
rect 583392 701752 583444 701758
rect 583392 701694 583444 701700
rect 583208 701616 583260 701622
rect 583208 701558 583260 701564
rect 583024 701480 583076 701486
rect 583024 701422 583076 701428
rect 582840 701344 582892 701350
rect 582840 701286 582892 701292
rect 582654 700360 582710 700369
rect 582654 700295 582710 700304
rect 582668 272241 582696 700295
rect 582852 312089 582880 701286
rect 582932 701276 582984 701282
rect 582932 701218 582984 701224
rect 582944 325281 582972 701218
rect 583036 365129 583064 701422
rect 583116 700256 583168 700262
rect 583116 700198 583168 700204
rect 583128 378457 583156 700198
rect 583220 418305 583248 701558
rect 583300 701548 583352 701554
rect 583300 701490 583352 701496
rect 583312 431633 583340 701490
rect 583404 484673 583432 701694
rect 583496 525065 583524 701898
rect 583576 701888 583628 701894
rect 583576 701830 583628 701836
rect 583588 538121 583616 701830
rect 583760 701208 583812 701214
rect 583760 701150 583812 701156
rect 583668 700324 583720 700330
rect 583668 700266 583720 700272
rect 583680 578241 583708 700266
rect 583666 578232 583722 578241
rect 583666 578167 583722 578176
rect 583574 538112 583630 538121
rect 583574 538047 583630 538056
rect 583482 525056 583538 525065
rect 583482 524991 583538 525000
rect 583390 484664 583446 484673
rect 583390 484599 583446 484608
rect 583298 431624 583354 431633
rect 583298 431559 583354 431568
rect 583206 418296 583262 418305
rect 583206 418231 583262 418240
rect 583114 378448 583170 378457
rect 583114 378383 583170 378392
rect 583022 365120 583078 365129
rect 583022 365055 583078 365064
rect 582930 325272 582986 325281
rect 582930 325207 582986 325216
rect 582838 312080 582894 312089
rect 582838 312015 582894 312024
rect 583772 299305 583800 701150
rect 583758 299296 583814 299305
rect 583758 299231 583814 299240
rect 582654 272232 582710 272241
rect 582654 272167 582710 272176
rect 582932 245608 582984 245614
rect 582930 245576 582932 245585
rect 582984 245576 582986 245585
rect 582930 245511 582986 245520
rect 582562 232384 582618 232393
rect 582562 232319 582618 232328
rect 582470 152688 582526 152697
rect 582470 152623 582526 152632
rect 582378 139360 582434 139369
rect 582378 139295 582434 139304
rect 582472 126064 582524 126070
rect 582470 126032 582472 126041
rect 582524 126032 582526 126041
rect 582470 125967 582526 125976
rect 580828 16546 580948 16574
rect 581196 16546 581776 16574
rect 580264 10396 580316 10402
rect 580264 10338 580316 10344
rect 580276 6633 580304 10338
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 580920 3482 580948 16546
rect 580920 3454 581040 3482
rect 578608 3052 578660 3058
rect 578608 2994 578660 3000
rect 579620 3052 579672 3058
rect 579620 2994 579672 3000
rect 578620 480 578648 2994
rect 581012 480 581040 3454
rect 581748 490 581776 16546
rect 583392 3528 583444 3534
rect 583392 3470 583444 3476
rect 582024 598 582236 626
rect 582024 490 582052 598
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 462 582052 490
rect 582208 480 582236 598
rect 583404 480 583432 3470
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3054 671200 3110 671256
rect 3330 619112 3386 619168
rect 3238 606056 3294 606112
rect 3238 462576 3294 462632
rect 3330 449520 3386 449576
rect 2962 410488 3018 410544
rect 3238 397432 3294 397488
rect 3514 658180 3516 658200
rect 3516 658180 3568 658200
rect 3568 658180 3570 658200
rect 3514 658144 3570 658180
rect 3514 633256 3570 633312
rect 3514 632032 3570 632088
rect 3514 580896 3570 580952
rect 3514 579944 3570 580000
rect 3514 566888 3570 566944
rect 3514 553832 3570 553888
rect 3514 514800 3570 514856
rect 3514 501744 3570 501800
rect 18602 701256 18658 701312
rect 3514 423580 3516 423600
rect 3516 423580 3568 423600
rect 3568 423580 3570 423600
rect 3514 423544 3570 423580
rect 21362 700712 21418 700768
rect 3514 371320 3570 371376
rect 3422 358400 3478 358456
rect 3146 345344 3202 345400
rect 3422 306176 3478 306232
rect 3054 293120 3110 293176
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 3422 202816 3478 202872
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3330 33088 3386 33144
rect 3330 32408 3386 32464
rect 3422 20576 3478 20632
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 29642 701120 29698 701176
rect 40498 700984 40554 701040
rect 32402 700032 32458 700088
rect 53194 699760 53250 699816
rect 68282 699896 68338 699952
rect 79322 701392 79378 701448
rect 105542 701528 105598 701584
rect 330666 703704 330722 703760
rect 165158 701800 165214 701856
rect 164514 701664 164570 701720
rect 164790 701664 164846 701720
rect 165342 701664 165398 701720
rect 194414 702072 194470 702128
rect 201314 701664 201370 701720
rect 212354 702208 212410 702264
rect 208812 701936 208868 701992
rect 205362 701800 205418 701856
rect 223394 702344 223450 702400
rect 227074 702344 227130 702400
rect 215850 701800 215906 701856
rect 218978 701800 219034 701856
rect 219622 701800 219678 701856
rect 226890 701800 226946 701856
rect 227074 701800 227130 701856
rect 234526 702344 234582 702400
rect 237930 702344 237986 702400
rect 264426 702344 264482 702400
rect 297546 702752 297602 702808
rect 286506 702616 286562 702672
rect 319626 703296 319682 703352
rect 315946 703160 316002 703216
rect 308586 702888 308642 702944
rect 300904 701936 300960 701992
rect 312266 702208 312322 702264
rect 326986 702208 327042 702264
rect 330206 702208 330262 702264
rect 334438 703840 334494 703896
rect 362498 703432 362554 703488
rect 350446 702480 350502 702536
rect 358726 702480 358782 702536
rect 361762 702480 361818 702536
rect 358726 702092 358782 702128
rect 358726 702072 358728 702092
rect 358728 702072 358780 702092
rect 358780 702072 358782 702092
rect 360290 702092 360346 702128
rect 360290 702072 360292 702092
rect 360292 702072 360344 702092
rect 360344 702072 360346 702092
rect 367190 702480 367246 702536
rect 418526 703568 418582 703624
rect 559378 703704 559434 703760
rect 429566 703024 429622 703080
rect 419354 702480 419410 702536
rect 481086 702480 481142 702536
rect 503258 702208 503314 702264
rect 510618 701528 510674 701584
rect 499670 701392 499726 701448
rect 488538 701256 488594 701312
rect 494794 701256 494850 701312
rect 506938 701256 506994 701312
rect 532698 702072 532754 702128
rect 514298 701120 514354 701176
rect 517978 701120 518034 701176
rect 521750 701120 521806 701176
rect 525430 701120 525486 701176
rect 527178 701120 527234 701176
rect 529018 701120 529074 701176
rect 536378 701120 536434 701176
rect 577042 703196 577044 703216
rect 577044 703196 577096 703216
rect 577096 703196 577098 703216
rect 577042 703160 577098 703196
rect 576950 702480 577006 702536
rect 582562 701800 582618 701856
rect 582470 701664 582526 701720
rect 573178 701120 573234 701176
rect 580538 701120 580594 701176
rect 582378 700168 582434 700224
rect 231214 280744 231270 280800
rect 233974 280880 234030 280936
rect 245014 280744 245070 280800
rect 580170 258848 580226 258904
rect 579986 219000 580042 219056
rect 580170 179152 580226 179208
rect 580170 112784 580226 112840
rect 579894 59608 579950 59664
rect 580446 86128 580502 86184
rect 580354 72936 580410 72992
rect 580262 46280 580318 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 582654 700304 582710 700360
rect 583666 578176 583722 578232
rect 583574 538056 583630 538112
rect 583482 525000 583538 525056
rect 583390 484608 583446 484664
rect 583298 431568 583354 431624
rect 583206 418240 583262 418296
rect 583114 378392 583170 378448
rect 583022 365064 583078 365120
rect 582930 325216 582986 325272
rect 582838 312024 582894 312080
rect 583758 299240 583814 299296
rect 582654 272176 582710 272232
rect 582930 245556 582932 245576
rect 582932 245556 582984 245576
rect 582984 245556 582986 245576
rect 582930 245520 582986 245556
rect 582562 232328 582618 232384
rect 582470 152632 582526 152688
rect 582378 139304 582434 139360
rect 582470 126012 582472 126032
rect 582472 126012 582524 126032
rect 582524 126012 582526 126032
rect 582470 125976 582526 126012
rect 580262 6568 580318 6624
<< metal3 >>
rect 334433 703898 334499 703901
rect 366950 703898 366956 703900
rect 334433 703896 366956 703898
rect 334433 703840 334438 703896
rect 334494 703840 366956 703896
rect 334433 703838 366956 703840
rect 334433 703835 334499 703838
rect 366950 703836 366956 703838
rect 367020 703836 367026 703900
rect 330661 703762 330727 703765
rect 559373 703762 559439 703765
rect 330661 703760 559439 703762
rect 330661 703704 330666 703760
rect 330722 703704 559378 703760
rect 559434 703704 559439 703760
rect 330661 703702 559439 703704
rect 330661 703699 330727 703702
rect 559373 703699 559439 703702
rect 324262 703564 324268 703628
rect 324332 703626 324338 703628
rect 418521 703626 418587 703629
rect 324332 703624 418587 703626
rect 324332 703568 418526 703624
rect 418582 703568 418587 703624
rect 324332 703566 418587 703568
rect 324332 703564 324338 703566
rect 418521 703563 418587 703566
rect 362493 703490 362559 703493
rect 580206 703490 580212 703492
rect 362493 703488 580212 703490
rect 362493 703432 362498 703488
rect 362554 703432 580212 703488
rect 362493 703430 580212 703432
rect 362493 703427 362559 703430
rect 580206 703428 580212 703430
rect 580276 703428 580282 703492
rect 319621 703354 319687 703357
rect 580022 703354 580028 703356
rect 319621 703352 580028 703354
rect 319621 703296 319626 703352
rect 319682 703296 580028 703352
rect 319621 703294 580028 703296
rect 319621 703291 319687 703294
rect 580022 703292 580028 703294
rect 580092 703292 580098 703356
rect 315941 703218 316007 703221
rect 577037 703218 577103 703221
rect 577262 703218 577268 703220
rect 315941 703216 567210 703218
rect 315941 703160 315946 703216
rect 316002 703160 567210 703216
rect 315941 703158 567210 703160
rect 315941 703155 316007 703158
rect 164918 703020 164924 703084
rect 164988 703082 164994 703084
rect 429561 703082 429627 703085
rect 164988 703080 429627 703082
rect 164988 703024 429566 703080
rect 429622 703024 429627 703080
rect 164988 703022 429627 703024
rect 567150 703082 567210 703158
rect 577037 703216 577268 703218
rect 577037 703160 577042 703216
rect 577098 703160 577268 703216
rect 577037 703158 577268 703160
rect 577037 703155 577103 703158
rect 577262 703156 577268 703158
rect 577332 703156 577338 703220
rect 577630 703082 577636 703084
rect 567150 703022 577636 703082
rect 164988 703020 164994 703022
rect 429561 703019 429627 703022
rect 577630 703020 577636 703022
rect 577700 703020 577706 703084
rect 308581 702946 308647 702949
rect 580758 702946 580764 702948
rect 308581 702944 580764 702946
rect 308581 702888 308586 702944
rect 308642 702888 580764 702944
rect 308581 702886 580764 702888
rect 308581 702883 308647 702886
rect 580758 702884 580764 702886
rect 580828 702884 580834 702948
rect 297541 702810 297607 702813
rect 580574 702810 580580 702812
rect 297541 702808 580580 702810
rect 297541 702752 297546 702808
rect 297602 702752 580580 702808
rect 297541 702750 580580 702752
rect 297541 702747 297607 702750
rect 580574 702748 580580 702750
rect 580644 702748 580650 702812
rect 286501 702674 286567 702677
rect 580390 702674 580396 702676
rect 286501 702672 580396 702674
rect 286501 702616 286506 702672
rect 286562 702616 580396 702672
rect 286501 702614 580396 702616
rect 286501 702611 286567 702614
rect 580390 702612 580396 702614
rect 580460 702612 580466 702676
rect 311750 702476 311756 702540
rect 311820 702538 311826 702540
rect 342846 702538 342852 702540
rect 311820 702478 342852 702538
rect 311820 702476 311826 702478
rect 342846 702476 342852 702478
rect 342916 702476 342922 702540
rect 350441 702538 350507 702541
rect 354622 702538 354628 702540
rect 350441 702536 354628 702538
rect 350441 702480 350446 702536
rect 350502 702480 354628 702536
rect 350441 702478 354628 702480
rect 350441 702475 350507 702478
rect 354622 702476 354628 702478
rect 354692 702476 354698 702540
rect 355174 702476 355180 702540
rect 355244 702538 355250 702540
rect 358721 702538 358787 702541
rect 355244 702536 358787 702538
rect 355244 702480 358726 702536
rect 358782 702480 358787 702536
rect 355244 702478 358787 702480
rect 355244 702476 355250 702478
rect 358721 702475 358787 702478
rect 360326 702476 360332 702540
rect 360396 702538 360402 702540
rect 361757 702538 361823 702541
rect 360396 702536 361823 702538
rect 360396 702480 361762 702536
rect 361818 702480 361823 702536
rect 360396 702478 361823 702480
rect 360396 702476 360402 702478
rect 361757 702475 361823 702478
rect 365662 702476 365668 702540
rect 365732 702538 365738 702540
rect 367185 702538 367251 702541
rect 419349 702540 419415 702541
rect 481081 702540 481147 702541
rect 419349 702538 419396 702540
rect 365732 702536 367251 702538
rect 365732 702480 367190 702536
rect 367246 702480 367251 702536
rect 365732 702478 367251 702480
rect 419304 702536 419396 702538
rect 419304 702480 419354 702536
rect 419304 702478 419396 702480
rect 365732 702476 365738 702478
rect 367185 702475 367251 702478
rect 419349 702476 419396 702478
rect 419460 702476 419466 702540
rect 481030 702538 481036 702540
rect 480990 702478 481036 702538
rect 481100 702536 481147 702540
rect 481142 702480 481147 702536
rect 481030 702476 481036 702478
rect 481100 702476 481147 702480
rect 419349 702475 419415 702476
rect 481081 702475 481147 702476
rect 576945 702538 577011 702541
rect 577078 702538 577084 702540
rect 576945 702536 577084 702538
rect 576945 702480 576950 702536
rect 577006 702480 577084 702536
rect 576945 702478 577084 702480
rect 576945 702475 577011 702478
rect 577078 702476 577084 702478
rect 577148 702476 577154 702540
rect 223389 702402 223455 702405
rect 227069 702402 227135 702405
rect 223389 702400 227135 702402
rect 223389 702344 223394 702400
rect 223450 702344 227074 702400
rect 227130 702344 227135 702400
rect 223389 702342 227135 702344
rect 223389 702339 223455 702342
rect 227069 702339 227135 702342
rect 234521 702402 234587 702405
rect 234654 702402 234660 702404
rect 234521 702400 234660 702402
rect 234521 702344 234526 702400
rect 234582 702344 234660 702400
rect 234521 702342 234660 702344
rect 234521 702339 234587 702342
rect 234654 702340 234660 702342
rect 234724 702340 234730 702404
rect 237414 702340 237420 702404
rect 237484 702402 237490 702404
rect 237925 702402 237991 702405
rect 237484 702400 237991 702402
rect 237484 702344 237930 702400
rect 237986 702344 237991 702400
rect 237484 702342 237991 702344
rect 237484 702340 237490 702342
rect 237925 702339 237991 702342
rect 264421 702402 264487 702405
rect 574686 702402 574692 702404
rect 264421 702400 574692 702402
rect 264421 702344 264426 702400
rect 264482 702344 574692 702400
rect 264421 702342 574692 702344
rect 264421 702339 264487 702342
rect 574686 702340 574692 702342
rect 574756 702340 574762 702404
rect 212349 702266 212415 702269
rect 312261 702268 312327 702269
rect 326981 702268 327047 702269
rect 244774 702266 244780 702268
rect 212349 702264 244780 702266
rect 212349 702208 212354 702264
rect 212410 702208 244780 702264
rect 212349 702206 244780 702208
rect 212349 702203 212415 702206
rect 244774 702204 244780 702206
rect 244844 702204 244850 702268
rect 312261 702264 312308 702268
rect 312372 702266 312378 702268
rect 312261 702208 312266 702264
rect 312261 702204 312308 702208
rect 312372 702206 312418 702266
rect 326981 702264 327028 702268
rect 327092 702266 327098 702268
rect 330201 702266 330267 702269
rect 503253 702266 503319 702269
rect 326981 702208 326986 702264
rect 312372 702204 312378 702206
rect 326981 702204 327028 702208
rect 327092 702206 327138 702266
rect 330201 702264 503319 702266
rect 330201 702208 330206 702264
rect 330262 702208 503258 702264
rect 503314 702208 503319 702264
rect 330201 702206 503319 702208
rect 327092 702204 327098 702206
rect 312261 702203 312327 702204
rect 326981 702203 327047 702204
rect 330201 702203 330267 702206
rect 503253 702203 503319 702206
rect 194409 702130 194475 702133
rect 357934 702130 357940 702132
rect 194409 702128 357940 702130
rect 194409 702072 194414 702128
rect 194470 702072 357940 702128
rect 194409 702070 357940 702072
rect 194409 702067 194475 702070
rect 357934 702068 357940 702070
rect 358004 702068 358010 702132
rect 358721 702130 358787 702133
rect 360142 702130 360148 702132
rect 358721 702128 360148 702130
rect 358721 702072 358726 702128
rect 358782 702072 360148 702128
rect 358721 702070 360148 702072
rect 358721 702067 358787 702070
rect 360142 702068 360148 702070
rect 360212 702068 360218 702132
rect 360285 702130 360351 702133
rect 532693 702130 532759 702133
rect 360285 702128 532759 702130
rect 360285 702072 360290 702128
rect 360346 702072 532698 702128
rect 532754 702072 532759 702128
rect 360285 702070 532759 702072
rect 360285 702067 360351 702070
rect 532693 702067 532759 702070
rect 208807 701994 208873 701997
rect 247718 701994 247724 701996
rect 208807 701992 247724 701994
rect 208807 701936 208812 701992
rect 208868 701936 247724 701992
rect 208807 701934 247724 701936
rect 208807 701931 208873 701934
rect 247718 701932 247724 701934
rect 247788 701932 247794 701996
rect 300899 701994 300965 701997
rect 575974 701994 575980 701996
rect 300899 701992 575980 701994
rect 300899 701936 300904 701992
rect 300960 701936 575980 701992
rect 300899 701934 575980 701936
rect 300899 701931 300965 701934
rect 575974 701932 575980 701934
rect 576044 701932 576050 701996
rect 165153 701860 165219 701861
rect 165102 701858 165108 701860
rect 165062 701798 165108 701858
rect 165172 701856 165219 701860
rect 165214 701800 165219 701856
rect 165102 701796 165108 701798
rect 165172 701796 165219 701800
rect 165153 701795 165219 701796
rect 205357 701860 205423 701861
rect 205357 701856 205404 701860
rect 205468 701858 205474 701860
rect 205357 701800 205362 701856
rect 205357 701796 205404 701800
rect 205468 701798 205514 701858
rect 205468 701796 205474 701798
rect 215334 701796 215340 701860
rect 215404 701858 215410 701860
rect 215845 701858 215911 701861
rect 218973 701860 219039 701861
rect 218973 701858 219020 701860
rect 215404 701856 215911 701858
rect 215404 701800 215850 701856
rect 215906 701800 215911 701856
rect 215404 701798 215911 701800
rect 218928 701856 219020 701858
rect 218928 701800 218978 701856
rect 218928 701798 219020 701800
rect 215404 701796 215410 701798
rect 205357 701795 205423 701796
rect 215845 701795 215911 701798
rect 218973 701796 219020 701798
rect 219084 701796 219090 701860
rect 219198 701796 219204 701860
rect 219268 701858 219274 701860
rect 219617 701858 219683 701861
rect 219268 701856 219683 701858
rect 219268 701800 219622 701856
rect 219678 701800 219683 701856
rect 219268 701798 219683 701800
rect 219268 701796 219274 701798
rect 218973 701795 219039 701796
rect 219617 701795 219683 701798
rect 226374 701796 226380 701860
rect 226444 701858 226450 701860
rect 226885 701858 226951 701861
rect 226444 701856 226951 701858
rect 226444 701800 226890 701856
rect 226946 701800 226951 701856
rect 226444 701798 226951 701800
rect 226444 701796 226450 701798
rect 226885 701795 226951 701798
rect 227069 701858 227135 701861
rect 582557 701858 582623 701861
rect 227069 701856 582623 701858
rect 227069 701800 227074 701856
rect 227130 701800 582562 701856
rect 582618 701800 582623 701856
rect 227069 701798 582623 701800
rect 227069 701795 227135 701798
rect 582557 701795 582623 701798
rect 164509 701724 164575 701725
rect 164785 701724 164851 701725
rect 165337 701724 165403 701725
rect 164509 701722 164556 701724
rect 164464 701720 164556 701722
rect 164464 701664 164514 701720
rect 164464 701662 164556 701664
rect 164509 701660 164556 701662
rect 164620 701660 164626 701724
rect 164734 701722 164740 701724
rect 164694 701662 164740 701722
rect 164804 701720 164851 701724
rect 165286 701722 165292 701724
rect 164846 701664 164851 701720
rect 164734 701660 164740 701662
rect 164804 701660 164851 701664
rect 165246 701662 165292 701722
rect 165356 701720 165403 701724
rect 165398 701664 165403 701720
rect 165286 701660 165292 701662
rect 165356 701660 165403 701664
rect 164509 701659 164575 701660
rect 164785 701659 164851 701660
rect 165337 701659 165403 701660
rect 201309 701722 201375 701725
rect 582465 701722 582531 701725
rect 201309 701720 582531 701722
rect 201309 701664 201314 701720
rect 201370 701664 582470 701720
rect 582526 701664 582531 701720
rect 201309 701662 582531 701664
rect 201309 701659 201375 701662
rect 582465 701659 582531 701662
rect 105537 701586 105603 701589
rect 510613 701586 510679 701589
rect 105537 701584 510679 701586
rect 105537 701528 105542 701584
rect 105598 701528 510618 701584
rect 510674 701528 510679 701584
rect 105537 701526 510679 701528
rect 105537 701523 105603 701526
rect 510613 701523 510679 701526
rect 79317 701450 79383 701453
rect 499665 701450 499731 701453
rect 79317 701448 499731 701450
rect 79317 701392 79322 701448
rect 79378 701392 499670 701448
rect 499726 701392 499731 701448
rect 79317 701390 499731 701392
rect 79317 701387 79383 701390
rect 499665 701387 499731 701390
rect 18597 701314 18663 701317
rect 488533 701314 488599 701317
rect 18597 701312 488599 701314
rect 18597 701256 18602 701312
rect 18658 701256 488538 701312
rect 488594 701256 488599 701312
rect 18597 701254 488599 701256
rect 18597 701251 18663 701254
rect 488533 701251 488599 701254
rect 494646 701252 494652 701316
rect 494716 701314 494722 701316
rect 494789 701314 494855 701317
rect 494716 701312 494855 701314
rect 494716 701256 494794 701312
rect 494850 701256 494855 701312
rect 494716 701254 494855 701256
rect 494716 701252 494722 701254
rect 494789 701251 494855 701254
rect 506422 701252 506428 701316
rect 506492 701314 506498 701316
rect 506933 701314 506999 701317
rect 506492 701312 506999 701314
rect 506492 701256 506938 701312
rect 506994 701256 506999 701312
rect 506492 701254 506999 701256
rect 506492 701252 506498 701254
rect 506933 701251 506999 701254
rect 29637 701178 29703 701181
rect 514293 701178 514359 701181
rect 29637 701176 514359 701178
rect 29637 701120 29642 701176
rect 29698 701120 514298 701176
rect 514354 701120 514359 701176
rect 29637 701118 514359 701120
rect 29637 701115 29703 701118
rect 514293 701115 514359 701118
rect 517646 701116 517652 701180
rect 517716 701178 517722 701180
rect 517973 701178 518039 701181
rect 521745 701180 521811 701181
rect 525425 701180 525491 701181
rect 521694 701178 521700 701180
rect 517716 701176 518039 701178
rect 517716 701120 517978 701176
rect 518034 701120 518039 701176
rect 517716 701118 518039 701120
rect 521654 701118 521700 701178
rect 521764 701176 521811 701180
rect 525374 701178 525380 701180
rect 521806 701120 521811 701176
rect 517716 701116 517722 701118
rect 517973 701115 518039 701118
rect 521694 701116 521700 701118
rect 521764 701116 521811 701120
rect 525334 701118 525380 701178
rect 525444 701176 525491 701180
rect 527173 701178 527239 701181
rect 525486 701120 525491 701176
rect 525374 701116 525380 701118
rect 525444 701116 525491 701120
rect 521745 701115 521811 701116
rect 525425 701115 525491 701116
rect 527038 701176 527239 701178
rect 527038 701120 527178 701176
rect 527234 701120 527239 701176
rect 527038 701118 527239 701120
rect 40493 701042 40559 701045
rect 324262 701042 324268 701044
rect 40493 701040 324268 701042
rect 40493 700984 40498 701040
rect 40554 700984 324268 701040
rect 40493 700982 324268 700984
rect 40493 700979 40559 700982
rect 324262 700980 324268 700982
rect 324332 700980 324338 701044
rect 342846 700980 342852 701044
rect 342916 701042 342922 701044
rect 355174 701042 355180 701044
rect 342916 700982 355180 701042
rect 342916 700980 342922 700982
rect 355174 700980 355180 700982
rect 355244 700980 355250 701044
rect 367502 700980 367508 701044
rect 367572 701042 367578 701044
rect 527038 701042 527098 701118
rect 527173 701115 527239 701118
rect 528318 701116 528324 701180
rect 528388 701178 528394 701180
rect 529013 701178 529079 701181
rect 528388 701176 529079 701178
rect 528388 701120 529018 701176
rect 529074 701120 529079 701176
rect 528388 701118 529079 701120
rect 528388 701116 528394 701118
rect 529013 701115 529079 701118
rect 533286 701116 533292 701180
rect 533356 701178 533362 701180
rect 536373 701178 536439 701181
rect 533356 701176 536439 701178
rect 533356 701120 536378 701176
rect 536434 701120 536439 701176
rect 533356 701118 536439 701120
rect 533356 701116 533362 701118
rect 536373 701115 536439 701118
rect 572662 701116 572668 701180
rect 572732 701178 572738 701180
rect 573173 701178 573239 701181
rect 572732 701176 573239 701178
rect 572732 701120 573178 701176
rect 573234 701120 573239 701176
rect 572732 701118 573239 701120
rect 572732 701116 572738 701118
rect 573173 701115 573239 701118
rect 577446 701116 577452 701180
rect 577516 701178 577522 701180
rect 580533 701178 580599 701181
rect 577516 701176 580599 701178
rect 577516 701120 580538 701176
rect 580594 701120 580599 701176
rect 577516 701118 580599 701120
rect 577516 701116 577522 701118
rect 580533 701115 580599 701118
rect 367572 700982 527098 701042
rect 367572 700980 367578 700982
rect 219014 700844 219020 700908
rect 219084 700906 219090 700908
rect 311750 700906 311756 700908
rect 219084 700846 311756 700906
rect 219084 700844 219090 700846
rect 311750 700844 311756 700846
rect 311820 700844 311826 700908
rect 354806 700844 354812 700908
rect 354876 700906 354882 700908
rect 494646 700906 494652 700908
rect 354876 700846 494652 700906
rect 354876 700844 354882 700846
rect 494646 700844 494652 700846
rect 494716 700844 494722 700908
rect 21357 700770 21423 700773
rect 365662 700770 365668 700772
rect 21357 700768 365668 700770
rect 21357 700712 21362 700768
rect 21418 700712 365668 700768
rect 21357 700710 365668 700712
rect 21357 700707 21423 700710
rect 365662 700708 365668 700710
rect 365732 700708 365738 700772
rect 419390 700708 419396 700772
rect 419460 700770 419466 700772
rect 579838 700770 579844 700772
rect 419460 700710 579844 700770
rect 419460 700708 419466 700710
rect 579838 700708 579844 700710
rect 579908 700708 579914 700772
rect 327022 700572 327028 700636
rect 327092 700634 327098 700636
rect 578734 700634 578740 700636
rect 327092 700574 578740 700634
rect 327092 700572 327098 700574
rect 578734 700572 578740 700574
rect 578804 700572 578810 700636
rect 312302 700436 312308 700500
rect 312372 700498 312378 700500
rect 574870 700498 574876 700500
rect 312372 700438 574876 700498
rect 312372 700436 312378 700438
rect 574870 700436 574876 700438
rect 574940 700436 574946 700500
rect 234654 700300 234660 700364
rect 234724 700362 234730 700364
rect 582649 700362 582715 700365
rect 234724 700360 582715 700362
rect 234724 700304 582654 700360
rect 582710 700304 582715 700360
rect 234724 700302 582715 700304
rect 234724 700300 234730 700302
rect 582649 700299 582715 700302
rect 205398 700164 205404 700228
rect 205468 700226 205474 700228
rect 582373 700226 582439 700229
rect 205468 700224 582439 700226
rect 205468 700168 582378 700224
rect 582434 700168 582439 700224
rect 205468 700166 582439 700168
rect 205468 700164 205474 700166
rect 582373 700163 582439 700166
rect 32397 700090 32463 700093
rect 481030 700090 481036 700092
rect 32397 700088 481036 700090
rect 32397 700032 32402 700088
rect 32458 700032 481036 700088
rect 32397 700030 481036 700032
rect 32397 700027 32463 700030
rect 481030 700028 481036 700030
rect 481100 700028 481106 700092
rect 68277 699954 68343 699957
rect 525374 699954 525380 699956
rect 68277 699952 525380 699954
rect 68277 699896 68282 699952
rect 68338 699896 525380 699952
rect 68277 699894 525380 699896
rect 68277 699891 68343 699894
rect 525374 699892 525380 699894
rect 525444 699892 525450 699956
rect 53189 699818 53255 699821
rect 521694 699818 521700 699820
rect 53189 699816 521700 699818
rect 53189 699760 53194 699816
rect 53250 699760 521700 699816
rect 53189 699758 521700 699760
rect 53189 699755 53255 699758
rect 521694 699756 521700 699758
rect 521764 699756 521770 699820
rect -960 697220 480 697460
rect 579838 697172 579844 697236
rect 579908 697234 579914 697236
rect 583520 697234 584960 697324
rect 579908 697174 584960 697234
rect 579908 697172 579914 697174
rect 583520 697084 584960 697174
rect 164918 684450 164924 684452
rect -960 684314 480 684404
rect 6870 684390 164924 684450
rect 6870 684314 6930 684390
rect 164918 684388 164924 684390
rect 164988 684388 164994 684452
rect -960 684254 6930 684314
rect -960 684164 480 684254
rect 578734 683844 578740 683908
rect 578804 683906 578810 683908
rect 583520 683906 584960 683996
rect 578804 683846 584960 683906
rect 578804 683844 578810 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3049 671258 3115 671261
rect -960 671256 3115 671258
rect -960 671200 3054 671256
rect 3110 671200 3115 671256
rect -960 671198 3115 671200
rect -960 671108 480 671198
rect 3049 671195 3115 671198
rect 580022 670652 580028 670716
rect 580092 670714 580098 670716
rect 583520 670714 584960 670804
rect 580092 670654 584960 670714
rect 580092 670652 580098 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 644058 584960 644148
rect 583342 643998 584960 644058
rect 583342 643922 583402 643998
rect 583520 643922 584960 643998
rect 583342 643908 584960 643922
rect 583342 643862 583586 643908
rect 574870 643180 574876 643244
rect 574940 643242 574946 643244
rect 583526 643242 583586 643862
rect 574940 643182 583586 643242
rect 574940 643180 574946 643182
rect 3509 633314 3575 633317
rect 164734 633314 164740 633316
rect 3509 633312 164740 633314
rect 3509 633256 3514 633312
rect 3570 633256 164740 633312
rect 3509 633254 164740 633256
rect 3509 633251 3575 633254
rect 164734 633252 164740 633254
rect 164804 633252 164810 633316
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 577630 630804 577636 630868
rect 577700 630866 577706 630868
rect 583520 630866 584960 630956
rect 577700 630806 584960 630866
rect 577700 630804 577706 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3325 619170 3391 619173
rect -960 619168 3391 619170
rect -960 619112 3330 619168
rect 3386 619112 3391 619168
rect -960 619110 3391 619112
rect -960 619020 480 619110
rect 3325 619107 3391 619110
rect 580758 617476 580764 617540
rect 580828 617538 580834 617540
rect 583520 617538 584960 617628
rect 580828 617478 584960 617538
rect 580828 617476 580834 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 575974 590956 575980 591020
rect 576044 591018 576050 591020
rect 583520 591018 584960 591108
rect 576044 590958 584960 591018
rect 576044 590956 576050 590958
rect 583520 590868 584960 590958
rect 3509 580954 3575 580957
rect 164550 580954 164556 580956
rect 3509 580952 164556 580954
rect 3509 580896 3514 580952
rect 3570 580896 164556 580952
rect 3509 580894 164556 580896
rect 3509 580891 3575 580894
rect 164550 580892 164556 580894
rect 164620 580892 164626 580956
rect -960 580002 480 580092
rect 3509 580002 3575 580005
rect -960 580000 3575 580002
rect -960 579944 3514 580000
rect 3570 579944 3575 580000
rect -960 579942 3575 579944
rect -960 579852 480 579942
rect 3509 579939 3575 579942
rect 583661 578234 583727 578237
rect 583526 578232 583727 578234
rect 583526 578176 583666 578232
rect 583722 578176 583727 578232
rect 583526 578174 583727 578176
rect 583526 577826 583586 578174
rect 583661 578171 583727 578174
rect 583342 577780 583586 577826
rect 583342 577766 584960 577780
rect 583342 577690 583402 577766
rect 583520 577690 584960 577766
rect 583342 577630 584960 577690
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 580574 564300 580580 564364
rect 580644 564362 580650 564364
rect 583520 564362 584960 564452
rect 580644 564302 584960 564362
rect 580644 564300 580650 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3509 553890 3575 553893
rect -960 553888 3575 553890
rect -960 553832 3514 553888
rect 3570 553832 3575 553888
rect -960 553830 3575 553832
rect -960 553740 480 553830
rect 3509 553827 3575 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583569 538114 583635 538117
rect 583526 538112 583635 538114
rect 583526 538056 583574 538112
rect 583630 538056 583635 538112
rect 583526 538051 583635 538056
rect 583526 537978 583586 538051
rect 583342 537932 583586 537978
rect 583342 537918 584960 537932
rect 583342 537842 583402 537918
rect 583520 537842 584960 537918
rect 583342 537782 584960 537842
rect 583520 537692 584960 537782
rect 165286 528458 165292 528460
rect 430 528398 165292 528458
rect 430 528186 490 528398
rect 165286 528396 165292 528398
rect 165356 528396 165362 528460
rect 430 528126 674 528186
rect -960 527914 480 528004
rect 614 527914 674 528126
rect -960 527854 674 527914
rect -960 527764 480 527854
rect 583477 525058 583543 525061
rect 583477 525056 583586 525058
rect 583477 525000 583482 525056
rect 583538 525000 583586 525056
rect 583477 524995 583586 525000
rect 583526 524650 583586 524995
rect 583342 524604 583586 524650
rect 583342 524590 584960 524604
rect 583342 524514 583402 524590
rect 583520 524514 584960 524590
rect 583342 524454 584960 524514
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580390 511260 580396 511324
rect 580460 511322 580466 511324
rect 583520 511322 584960 511412
rect 580460 511262 584960 511322
rect 580460 511260 580466 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583385 484666 583451 484669
rect 583520 484666 584960 484756
rect 583385 484664 584960 484666
rect 583385 484608 583390 484664
rect 583446 484608 584960 484664
rect 583385 484606 584960 484608
rect 583385 484603 583451 484606
rect 583520 484516 584960 484606
rect 165102 476098 165108 476100
rect 6870 476038 165108 476098
rect -960 475690 480 475780
rect 6870 475690 6930 476038
rect 165102 476036 165108 476038
rect 165172 476036 165178 476100
rect -960 475630 6930 475690
rect -960 475540 480 475630
rect 577078 471412 577084 471476
rect 577148 471474 577154 471476
rect 583520 471474 584960 471564
rect 577148 471414 584960 471474
rect 577148 471412 577154 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580206 458084 580212 458148
rect 580276 458146 580282 458148
rect 583520 458146 584960 458236
rect 580276 458086 584960 458146
rect 580276 458084 580282 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583293 431626 583359 431629
rect 583520 431626 584960 431716
rect 583293 431624 584960 431626
rect 583293 431568 583298 431624
rect 583354 431568 584960 431624
rect 583293 431566 584960 431568
rect 583293 431563 583359 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 583201 418298 583267 418301
rect 583520 418298 584960 418388
rect 583201 418296 584960 418298
rect 583201 418240 583206 418296
rect 583262 418240 584960 418296
rect 583201 418238 584960 418240
rect 583201 418235 583267 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 583520 404970 584960 405060
rect 583342 404910 584960 404970
rect 583342 404834 583402 404910
rect 583520 404834 584960 404910
rect 583342 404820 584960 404834
rect 583342 404774 583586 404820
rect 574686 404364 574692 404428
rect 574756 404426 574762 404428
rect 583526 404426 583586 404774
rect 574756 404366 583586 404426
rect 574756 404364 574762 404366
rect -960 397490 480 397580
rect 3233 397490 3299 397493
rect -960 397488 3299 397490
rect -960 397432 3238 397488
rect 3294 397432 3299 397488
rect -960 397430 3299 397432
rect -960 397340 480 397430
rect 3233 397427 3299 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583109 378450 583175 378453
rect 583520 378450 584960 378540
rect 583109 378448 584960 378450
rect 583109 378392 583114 378448
rect 583170 378392 584960 378448
rect 583109 378390 584960 378392
rect 583109 378387 583175 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 583017 365122 583083 365125
rect 583520 365122 584960 365212
rect 583017 365120 584960 365122
rect 583017 365064 583022 365120
rect 583078 365064 584960 365120
rect 583017 365062 584960 365064
rect 583017 365059 583083 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 577262 351868 577268 351932
rect 577332 351930 577338 351932
rect 583520 351930 584960 352020
rect 577332 351870 584960 351930
rect 577332 351868 577338 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 582925 325274 582991 325277
rect 583520 325274 584960 325364
rect 582925 325272 584960 325274
rect 582925 325216 582930 325272
rect 582986 325216 584960 325272
rect 582925 325214 584960 325216
rect 582925 325211 582991 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect -960 319230 6930 319290
rect -960 319140 480 319230
rect 6870 318882 6930 319230
rect 164734 318882 164740 318884
rect 6870 318822 164740 318882
rect 164734 318820 164740 318822
rect 164804 318820 164810 318884
rect 582833 312082 582899 312085
rect 583520 312082 584960 312172
rect 582833 312080 584960 312082
rect 582833 312024 582838 312080
rect 582894 312024 584960 312080
rect 582833 312022 584960 312024
rect 582833 312019 582899 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 583753 299298 583819 299301
rect 583710 299296 583819 299298
rect 583710 299240 583758 299296
rect 583814 299240 583819 299296
rect 583710 299235 583819 299240
rect 583710 298890 583770 299235
rect 583342 298844 583770 298890
rect 583342 298830 584960 298844
rect 583342 298754 583402 298830
rect 583520 298754 584960 298830
rect 583342 298694 584960 298754
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 583520 285276 584960 285516
rect 164734 283732 164740 283796
rect 164804 283794 164810 283796
rect 506422 283794 506428 283796
rect 164804 283734 506428 283794
rect 164804 283732 164810 283734
rect 506422 283732 506428 283734
rect 506492 283732 506498 283796
rect 226374 280876 226380 280940
rect 226444 280938 226450 280940
rect 233969 280938 234035 280941
rect 226444 280936 234035 280938
rect 226444 280880 233974 280936
rect 234030 280880 234035 280936
rect 226444 280878 234035 280880
rect 226444 280876 226450 280878
rect 233969 280875 234035 280878
rect 215334 280740 215340 280804
rect 215404 280802 215410 280804
rect 231209 280802 231275 280805
rect 215404 280800 231275 280802
rect 215404 280744 231214 280800
rect 231270 280744 231275 280800
rect 215404 280742 231275 280744
rect 215404 280740 215410 280742
rect 231209 280739 231275 280742
rect 237414 280740 237420 280804
rect 237484 280802 237490 280804
rect 245009 280802 245075 280805
rect 237484 280800 245075 280802
rect 237484 280744 245014 280800
rect 245070 280744 245075 280800
rect 237484 280742 245075 280744
rect 237484 280740 237490 280742
rect 245009 280739 245075 280742
rect -960 279972 480 280212
rect 582649 272234 582715 272237
rect 583520 272234 584960 272324
rect 582649 272232 584960 272234
rect 582649 272176 582654 272232
rect 582710 272176 584960 272232
rect 582649 272174 584960 272176
rect 582649 272171 582715 272174
rect 583520 272084 584960 272174
rect 517830 267746 517836 267748
rect 430 267686 517836 267746
rect 430 267474 490 267686
rect 517830 267684 517836 267686
rect 517900 267684 517906 267748
rect 430 267414 674 267474
rect -960 267202 480 267292
rect 614 267202 674 267414
rect -960 267142 674 267202
rect -960 267052 480 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 582925 245578 582991 245581
rect 583520 245578 584960 245668
rect 582925 245576 584960 245578
rect 582925 245520 582930 245576
rect 582986 245520 584960 245576
rect 582925 245518 584960 245520
rect 582925 245515 582991 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 582557 232386 582623 232389
rect 583520 232386 584960 232476
rect 582557 232384 584960 232386
rect 582557 232328 582562 232384
rect 582618 232328 584960 232384
rect 582557 232326 584960 232328
rect 582557 232323 582623 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579981 219058 580047 219061
rect 583520 219058 584960 219148
rect 579981 219056 584960 219058
rect 579981 219000 579986 219056
rect 580042 219000 584960 219056
rect 579981 218998 584960 219000
rect 579981 218995 580047 218998
rect 583520 218908 584960 218998
rect 528318 215250 528324 215252
rect 6870 215190 528324 215250
rect -960 214978 480 215068
rect 6870 214978 6930 215190
rect 528318 215188 528324 215190
rect 528388 215188 528394 215252
rect -960 214918 6930 214978
rect -960 214828 480 214918
rect 219382 205668 219388 205732
rect 219452 205730 219458 205732
rect 583520 205730 584960 205820
rect 219452 205670 584960 205730
rect 219452 205668 219458 205670
rect 583520 205580 584960 205670
rect 3417 202874 3483 202877
rect 533286 202874 533292 202876
rect 3417 202872 533292 202874
rect 3417 202816 3422 202872
rect 3478 202816 533292 202872
rect 3417 202814 533292 202816
rect 3417 202811 3483 202814
rect 533286 202812 533292 202814
rect 533356 202812 533362 202876
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 583520 192538 584960 192628
rect 583342 192478 584960 192538
rect 583342 192402 583402 192478
rect 583520 192402 584960 192478
rect 583342 192388 584960 192402
rect 583342 192342 583586 192388
rect 244774 191796 244780 191860
rect 244844 191858 244850 191860
rect 583526 191858 583586 192342
rect 244844 191798 583586 191858
rect 244844 191796 244850 191798
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 583520 165882 584960 165972
rect 567150 165822 584960 165882
rect 247718 165684 247724 165748
rect 247788 165746 247794 165748
rect 567150 165746 567210 165822
rect 247788 165686 567210 165746
rect 583520 165732 584960 165822
rect 247788 165684 247794 165686
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 582465 152690 582531 152693
rect 583520 152690 584960 152780
rect 582465 152688 584960 152690
rect 582465 152632 582470 152688
rect 582526 152632 584960 152688
rect 582465 152630 584960 152632
rect 582465 152627 582531 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 582373 139362 582439 139365
rect 583520 139362 584960 139452
rect 582373 139360 584960 139362
rect 582373 139304 582378 139360
rect 582434 139304 584960 139360
rect 582373 139302 584960 139304
rect 582373 139299 582439 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 582465 126034 582531 126037
rect 583520 126034 584960 126124
rect 582465 126032 584960 126034
rect 582465 125976 582470 126032
rect 582526 125976 584960 126032
rect 582465 125974 584960 125976
rect 582465 125971 582531 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 357934 99452 357940 99516
rect 358004 99514 358010 99516
rect 583520 99514 584960 99604
rect 358004 99454 584960 99514
rect 358004 99452 358010 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 580441 86186 580507 86189
rect 583520 86186 584960 86276
rect 580441 86184 584960 86186
rect 580441 86128 580446 86184
rect 580502 86128 584960 86184
rect 580441 86126 584960 86128
rect 580441 86123 580507 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 579889 59666 579955 59669
rect 583520 59666 584960 59756
rect 579889 59664 584960 59666
rect 579889 59608 579894 59664
rect 579950 59608 584960 59664
rect 579889 59606 584960 59608
rect 579889 59603 579955 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580257 46338 580323 46341
rect 583520 46338 584960 46428
rect 580257 46336 584960 46338
rect 580257 46280 580262 46336
rect 580318 46280 584960 46336
rect 580257 46278 584960 46280
rect 580257 46275 580323 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 3325 33146 3391 33149
rect 572662 33146 572668 33148
rect 3325 33144 572668 33146
rect 3325 33088 3330 33144
rect 3386 33088 572668 33144
rect 3325 33086 572668 33088
rect 3325 33083 3391 33086
rect 572662 33084 572668 33086
rect 572732 33084 572738 33148
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3325 32466 3391 32469
rect -960 32464 3391 32466
rect -960 32408 3330 32464
rect 3386 32408 3391 32464
rect -960 32406 3391 32408
rect -960 32316 480 32406
rect 3325 32403 3391 32406
rect 3417 20634 3483 20637
rect 577446 20634 577452 20636
rect 3417 20632 577452 20634
rect 3417 20576 3422 20632
rect 3478 20576 577452 20632
rect 3417 20574 577452 20576
rect 3417 20571 3483 20574
rect 577446 20572 577452 20574
rect 577516 20572 577522 20636
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 366956 703836 367020 703900
rect 324268 703564 324332 703628
rect 580212 703428 580276 703492
rect 580028 703292 580092 703356
rect 164924 703020 164988 703084
rect 577268 703156 577332 703220
rect 577636 703020 577700 703084
rect 580764 702884 580828 702948
rect 580580 702748 580644 702812
rect 580396 702612 580460 702676
rect 311756 702476 311820 702540
rect 342852 702476 342916 702540
rect 354628 702476 354692 702540
rect 355180 702476 355244 702540
rect 360332 702476 360396 702540
rect 365668 702476 365732 702540
rect 419396 702536 419460 702540
rect 419396 702480 419410 702536
rect 419410 702480 419460 702536
rect 419396 702476 419460 702480
rect 481036 702536 481100 702540
rect 481036 702480 481086 702536
rect 481086 702480 481100 702536
rect 481036 702476 481100 702480
rect 577084 702476 577148 702540
rect 234660 702340 234724 702404
rect 237420 702340 237484 702404
rect 574692 702340 574756 702404
rect 244780 702204 244844 702268
rect 312308 702264 312372 702268
rect 312308 702208 312322 702264
rect 312322 702208 312372 702264
rect 312308 702204 312372 702208
rect 327028 702264 327092 702268
rect 327028 702208 327042 702264
rect 327042 702208 327092 702264
rect 327028 702204 327092 702208
rect 357940 702068 358004 702132
rect 360148 702068 360212 702132
rect 247724 701932 247788 701996
rect 575980 701932 576044 701996
rect 165108 701856 165172 701860
rect 165108 701800 165158 701856
rect 165158 701800 165172 701856
rect 165108 701796 165172 701800
rect 205404 701856 205468 701860
rect 205404 701800 205418 701856
rect 205418 701800 205468 701856
rect 205404 701796 205468 701800
rect 215340 701796 215404 701860
rect 219020 701856 219084 701860
rect 219020 701800 219034 701856
rect 219034 701800 219084 701856
rect 219020 701796 219084 701800
rect 219204 701796 219268 701860
rect 226380 701796 226444 701860
rect 164556 701720 164620 701724
rect 164556 701664 164570 701720
rect 164570 701664 164620 701720
rect 164556 701660 164620 701664
rect 164740 701720 164804 701724
rect 164740 701664 164790 701720
rect 164790 701664 164804 701720
rect 164740 701660 164804 701664
rect 165292 701720 165356 701724
rect 165292 701664 165342 701720
rect 165342 701664 165356 701720
rect 165292 701660 165356 701664
rect 494652 701252 494716 701316
rect 506428 701252 506492 701316
rect 517652 701116 517716 701180
rect 521700 701176 521764 701180
rect 521700 701120 521750 701176
rect 521750 701120 521764 701176
rect 521700 701116 521764 701120
rect 525380 701176 525444 701180
rect 525380 701120 525430 701176
rect 525430 701120 525444 701176
rect 525380 701116 525444 701120
rect 324268 700980 324332 701044
rect 342852 700980 342916 701044
rect 355180 700980 355244 701044
rect 367508 700980 367572 701044
rect 528324 701116 528388 701180
rect 533292 701116 533356 701180
rect 572668 701116 572732 701180
rect 577452 701116 577516 701180
rect 219020 700844 219084 700908
rect 311756 700844 311820 700908
rect 354812 700844 354876 700908
rect 494652 700844 494716 700908
rect 365668 700708 365732 700772
rect 419396 700708 419460 700772
rect 579844 700708 579908 700772
rect 327028 700572 327092 700636
rect 578740 700572 578804 700636
rect 312308 700436 312372 700500
rect 574876 700436 574940 700500
rect 234660 700300 234724 700364
rect 205404 700164 205468 700228
rect 481036 700028 481100 700092
rect 525380 699892 525444 699956
rect 521700 699756 521764 699820
rect 579844 697172 579908 697236
rect 164924 684388 164988 684452
rect 578740 683844 578804 683908
rect 580028 670652 580092 670716
rect 574876 643180 574940 643244
rect 164740 633252 164804 633316
rect 577636 630804 577700 630868
rect 580764 617476 580828 617540
rect 575980 590956 576044 591020
rect 164556 580892 164620 580956
rect 580580 564300 580644 564364
rect 165292 528396 165356 528460
rect 580396 511260 580460 511324
rect 165108 476036 165172 476100
rect 577084 471412 577148 471476
rect 580212 458084 580276 458148
rect 574692 404364 574756 404428
rect 577268 351868 577332 351932
rect 164740 318820 164804 318884
rect 164740 283732 164804 283796
rect 506428 283732 506492 283796
rect 226380 280876 226444 280940
rect 215340 280740 215404 280804
rect 237420 280740 237484 280804
rect 517836 267684 517900 267748
rect 528324 215188 528388 215252
rect 219388 205668 219452 205732
rect 533292 202812 533356 202876
rect 244780 191796 244844 191860
rect 247724 165684 247788 165748
rect 357940 99452 358004 99516
rect 572668 33084 572732 33148
rect 577452 20572 577516 20636
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 701792 164414 705242
rect 167514 703792 168134 707162
rect 171234 703792 171854 709082
rect 174954 703792 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 164923 703084 164989 703085
rect 164923 703020 164924 703084
rect 164988 703020 164989 703084
rect 164923 703019 164989 703020
rect 164555 701724 164621 701725
rect 164555 701660 164556 701724
rect 164620 701660 164621 701724
rect 164555 701659 164621 701660
rect 164739 701724 164805 701725
rect 164739 701660 164740 701724
rect 164804 701660 164805 701724
rect 164739 701659 164805 701660
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 164558 580957 164618 701659
rect 164742 633317 164802 701659
rect 164926 684453 164986 703019
rect 165107 701860 165173 701861
rect 165107 701796 165108 701860
rect 165172 701796 165173 701860
rect 165107 701795 165173 701796
rect 164923 684452 164989 684453
rect 164923 684388 164924 684452
rect 164988 684388 164989 684452
rect 164923 684387 164989 684388
rect 164739 633316 164805 633317
rect 164739 633252 164740 633316
rect 164804 633252 164805 633316
rect 164739 633251 164805 633252
rect 164555 580956 164621 580957
rect 164555 580892 164556 580956
rect 164620 580892 164621 580956
rect 164555 580891 164621 580892
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 165110 476101 165170 701795
rect 181794 701792 182414 704282
rect 185514 703792 186134 706202
rect 189234 703792 189854 708122
rect 192954 703792 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 701792 200414 705242
rect 203514 703792 204134 707162
rect 207234 703792 207854 709082
rect 210954 703792 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 205403 701860 205469 701861
rect 205403 701796 205404 701860
rect 205468 701796 205469 701860
rect 205403 701795 205469 701796
rect 215339 701860 215405 701861
rect 215339 701796 215340 701860
rect 215404 701796 215405 701860
rect 215339 701795 215405 701796
rect 165291 701724 165357 701725
rect 165291 701660 165292 701724
rect 165356 701660 165357 701724
rect 165291 701659 165357 701660
rect 165294 528461 165354 701659
rect 205406 700229 205466 701795
rect 205403 700228 205469 700229
rect 205403 700164 205404 700228
rect 205468 700164 205469 700228
rect 205403 700163 205469 700164
rect 167000 687454 167320 687486
rect 167000 687218 167042 687454
rect 167278 687218 167320 687454
rect 167000 687134 167320 687218
rect 167000 686898 167042 687134
rect 167278 686898 167320 687134
rect 167000 686866 167320 686898
rect 197720 687454 198040 687486
rect 197720 687218 197762 687454
rect 197998 687218 198040 687454
rect 197720 687134 198040 687218
rect 197720 686898 197762 687134
rect 197998 686898 198040 687134
rect 197720 686866 198040 686898
rect 182360 669454 182680 669486
rect 182360 669218 182402 669454
rect 182638 669218 182680 669454
rect 182360 669134 182680 669218
rect 182360 668898 182402 669134
rect 182638 668898 182680 669134
rect 182360 668866 182680 668898
rect 213080 669454 213400 669486
rect 213080 669218 213122 669454
rect 213358 669218 213400 669454
rect 213080 669134 213400 669218
rect 213080 668898 213122 669134
rect 213358 668898 213400 669134
rect 213080 668866 213400 668898
rect 167000 651454 167320 651486
rect 167000 651218 167042 651454
rect 167278 651218 167320 651454
rect 167000 651134 167320 651218
rect 167000 650898 167042 651134
rect 167278 650898 167320 651134
rect 167000 650866 167320 650898
rect 197720 651454 198040 651486
rect 197720 651218 197762 651454
rect 197998 651218 198040 651454
rect 197720 651134 198040 651218
rect 197720 650898 197762 651134
rect 197998 650898 198040 651134
rect 197720 650866 198040 650898
rect 182360 633454 182680 633486
rect 182360 633218 182402 633454
rect 182638 633218 182680 633454
rect 182360 633134 182680 633218
rect 182360 632898 182402 633134
rect 182638 632898 182680 633134
rect 182360 632866 182680 632898
rect 213080 633454 213400 633486
rect 213080 633218 213122 633454
rect 213358 633218 213400 633454
rect 213080 633134 213400 633218
rect 213080 632898 213122 633134
rect 213358 632898 213400 633134
rect 213080 632866 213400 632898
rect 167000 615454 167320 615486
rect 167000 615218 167042 615454
rect 167278 615218 167320 615454
rect 167000 615134 167320 615218
rect 167000 614898 167042 615134
rect 167278 614898 167320 615134
rect 167000 614866 167320 614898
rect 197720 615454 198040 615486
rect 197720 615218 197762 615454
rect 197998 615218 198040 615454
rect 197720 615134 198040 615218
rect 197720 614898 197762 615134
rect 197998 614898 198040 615134
rect 197720 614866 198040 614898
rect 182360 597454 182680 597486
rect 182360 597218 182402 597454
rect 182638 597218 182680 597454
rect 182360 597134 182680 597218
rect 182360 596898 182402 597134
rect 182638 596898 182680 597134
rect 182360 596866 182680 596898
rect 213080 597454 213400 597486
rect 213080 597218 213122 597454
rect 213358 597218 213400 597454
rect 213080 597134 213400 597218
rect 213080 596898 213122 597134
rect 213358 596898 213400 597134
rect 213080 596866 213400 596898
rect 167000 579454 167320 579486
rect 167000 579218 167042 579454
rect 167278 579218 167320 579454
rect 167000 579134 167320 579218
rect 167000 578898 167042 579134
rect 167278 578898 167320 579134
rect 167000 578866 167320 578898
rect 197720 579454 198040 579486
rect 197720 579218 197762 579454
rect 197998 579218 198040 579454
rect 197720 579134 198040 579218
rect 197720 578898 197762 579134
rect 197998 578898 198040 579134
rect 197720 578866 198040 578898
rect 182360 561454 182680 561486
rect 182360 561218 182402 561454
rect 182638 561218 182680 561454
rect 182360 561134 182680 561218
rect 182360 560898 182402 561134
rect 182638 560898 182680 561134
rect 182360 560866 182680 560898
rect 213080 561454 213400 561486
rect 213080 561218 213122 561454
rect 213358 561218 213400 561454
rect 213080 561134 213400 561218
rect 213080 560898 213122 561134
rect 213358 560898 213400 561134
rect 213080 560866 213400 560898
rect 167000 543454 167320 543486
rect 167000 543218 167042 543454
rect 167278 543218 167320 543454
rect 167000 543134 167320 543218
rect 167000 542898 167042 543134
rect 167278 542898 167320 543134
rect 167000 542866 167320 542898
rect 197720 543454 198040 543486
rect 197720 543218 197762 543454
rect 197998 543218 198040 543454
rect 197720 543134 198040 543218
rect 197720 542898 197762 543134
rect 197998 542898 198040 543134
rect 197720 542866 198040 542898
rect 165291 528460 165357 528461
rect 165291 528396 165292 528460
rect 165356 528396 165357 528460
rect 165291 528395 165357 528396
rect 182360 525454 182680 525486
rect 182360 525218 182402 525454
rect 182638 525218 182680 525454
rect 182360 525134 182680 525218
rect 182360 524898 182402 525134
rect 182638 524898 182680 525134
rect 182360 524866 182680 524898
rect 213080 525454 213400 525486
rect 213080 525218 213122 525454
rect 213358 525218 213400 525454
rect 213080 525134 213400 525218
rect 213080 524898 213122 525134
rect 213358 524898 213400 525134
rect 213080 524866 213400 524898
rect 167000 507454 167320 507486
rect 167000 507218 167042 507454
rect 167278 507218 167320 507454
rect 167000 507134 167320 507218
rect 167000 506898 167042 507134
rect 167278 506898 167320 507134
rect 167000 506866 167320 506898
rect 197720 507454 198040 507486
rect 197720 507218 197762 507454
rect 197998 507218 198040 507454
rect 197720 507134 198040 507218
rect 197720 506898 197762 507134
rect 197998 506898 198040 507134
rect 197720 506866 198040 506898
rect 182360 489454 182680 489486
rect 182360 489218 182402 489454
rect 182638 489218 182680 489454
rect 182360 489134 182680 489218
rect 182360 488898 182402 489134
rect 182638 488898 182680 489134
rect 182360 488866 182680 488898
rect 213080 489454 213400 489486
rect 213080 489218 213122 489454
rect 213358 489218 213400 489454
rect 213080 489134 213400 489218
rect 213080 488898 213122 489134
rect 213358 488898 213400 489134
rect 213080 488866 213400 488898
rect 165107 476100 165173 476101
rect 165107 476036 165108 476100
rect 165172 476036 165173 476100
rect 165107 476035 165173 476036
rect 167000 471454 167320 471486
rect 167000 471218 167042 471454
rect 167278 471218 167320 471454
rect 167000 471134 167320 471218
rect 167000 470898 167042 471134
rect 167278 470898 167320 471134
rect 167000 470866 167320 470898
rect 197720 471454 198040 471486
rect 197720 471218 197762 471454
rect 197998 471218 198040 471454
rect 197720 471134 198040 471218
rect 197720 470898 197762 471134
rect 197998 470898 198040 471134
rect 197720 470866 198040 470898
rect 182360 453454 182680 453486
rect 182360 453218 182402 453454
rect 182638 453218 182680 453454
rect 182360 453134 182680 453218
rect 182360 452898 182402 453134
rect 182638 452898 182680 453134
rect 182360 452866 182680 452898
rect 213080 453454 213400 453486
rect 213080 453218 213122 453454
rect 213358 453218 213400 453454
rect 213080 453134 213400 453218
rect 213080 452898 213122 453134
rect 213358 452898 213400 453134
rect 213080 452866 213400 452898
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 167000 435454 167320 435486
rect 167000 435218 167042 435454
rect 167278 435218 167320 435454
rect 167000 435134 167320 435218
rect 167000 434898 167042 435134
rect 167278 434898 167320 435134
rect 167000 434866 167320 434898
rect 197720 435454 198040 435486
rect 197720 435218 197762 435454
rect 197998 435218 198040 435454
rect 197720 435134 198040 435218
rect 197720 434898 197762 435134
rect 197998 434898 198040 435134
rect 197720 434866 198040 434898
rect 182360 417454 182680 417486
rect 182360 417218 182402 417454
rect 182638 417218 182680 417454
rect 182360 417134 182680 417218
rect 182360 416898 182402 417134
rect 182638 416898 182680 417134
rect 182360 416866 182680 416898
rect 213080 417454 213400 417486
rect 213080 417218 213122 417454
rect 213358 417218 213400 417454
rect 213080 417134 213400 417218
rect 213080 416898 213122 417134
rect 213358 416898 213400 417134
rect 213080 416866 213400 416898
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 167000 399454 167320 399486
rect 167000 399218 167042 399454
rect 167278 399218 167320 399454
rect 167000 399134 167320 399218
rect 167000 398898 167042 399134
rect 167278 398898 167320 399134
rect 167000 398866 167320 398898
rect 197720 399454 198040 399486
rect 197720 399218 197762 399454
rect 197998 399218 198040 399454
rect 197720 399134 198040 399218
rect 197720 398898 197762 399134
rect 197998 398898 198040 399134
rect 197720 398866 198040 398898
rect 182360 381454 182680 381486
rect 182360 381218 182402 381454
rect 182638 381218 182680 381454
rect 182360 381134 182680 381218
rect 182360 380898 182402 381134
rect 182638 380898 182680 381134
rect 182360 380866 182680 380898
rect 213080 381454 213400 381486
rect 213080 381218 213122 381454
rect 213358 381218 213400 381454
rect 213080 381134 213400 381218
rect 213080 380898 213122 381134
rect 213358 380898 213400 381134
rect 213080 380866 213400 380898
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 167000 363454 167320 363486
rect 167000 363218 167042 363454
rect 167278 363218 167320 363454
rect 167000 363134 167320 363218
rect 167000 362898 167042 363134
rect 167278 362898 167320 363134
rect 167000 362866 167320 362898
rect 197720 363454 198040 363486
rect 197720 363218 197762 363454
rect 197998 363218 198040 363454
rect 197720 363134 198040 363218
rect 197720 362898 197762 363134
rect 197998 362898 198040 363134
rect 197720 362866 198040 362898
rect 182360 345454 182680 345486
rect 182360 345218 182402 345454
rect 182638 345218 182680 345454
rect 182360 345134 182680 345218
rect 182360 344898 182402 345134
rect 182638 344898 182680 345134
rect 182360 344866 182680 344898
rect 213080 345454 213400 345486
rect 213080 345218 213122 345454
rect 213358 345218 213400 345454
rect 213080 345134 213400 345218
rect 213080 344898 213122 345134
rect 213358 344898 213400 345134
rect 213080 344866 213400 344898
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 167000 327454 167320 327486
rect 167000 327218 167042 327454
rect 167278 327218 167320 327454
rect 167000 327134 167320 327218
rect 167000 326898 167042 327134
rect 167278 326898 167320 327134
rect 167000 326866 167320 326898
rect 197720 327454 198040 327486
rect 197720 327218 197762 327454
rect 197998 327218 198040 327454
rect 197720 327134 198040 327218
rect 197720 326898 197762 327134
rect 197998 326898 198040 327134
rect 197720 326866 198040 326898
rect 164739 318884 164805 318885
rect 164739 318820 164740 318884
rect 164804 318820 164805 318884
rect 164739 318819 164805 318820
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 164742 283797 164802 318819
rect 182360 309454 182680 309486
rect 182360 309218 182402 309454
rect 182638 309218 182680 309454
rect 182360 309134 182680 309218
rect 182360 308898 182402 309134
rect 182638 308898 182680 309134
rect 182360 308866 182680 308898
rect 213080 309454 213400 309486
rect 213080 309218 213122 309454
rect 213358 309218 213400 309454
rect 213080 309134 213400 309218
rect 213080 308898 213122 309134
rect 213358 308898 213400 309134
rect 213080 308866 213400 308898
rect 167000 291454 167320 291486
rect 167000 291218 167042 291454
rect 167278 291218 167320 291454
rect 167000 291134 167320 291218
rect 167000 290898 167042 291134
rect 167278 290898 167320 291134
rect 167000 290866 167320 290898
rect 197720 291454 198040 291486
rect 197720 291218 197762 291454
rect 197998 291218 198040 291454
rect 197720 291134 198040 291218
rect 197720 290898 197762 291134
rect 197998 290898 198040 291134
rect 197720 290866 198040 290898
rect 164739 283796 164805 283797
rect 164739 283732 164740 283796
rect 164804 283732 164805 283796
rect 164739 283731 164805 283732
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 273454 164414 281792
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 277174 168134 279792
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 244894 171854 279792
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 248614 175574 279792
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 255454 182414 281792
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 259174 186134 279792
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 262894 189854 279792
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 266614 193574 279792
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 273454 200414 281792
rect 215342 280805 215402 701795
rect 217794 701792 218414 704282
rect 221514 703792 222134 706202
rect 225234 703792 225854 708122
rect 228954 703792 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 234659 702404 234725 702405
rect 234659 702340 234660 702404
rect 234724 702340 234725 702404
rect 234659 702339 234725 702340
rect 219019 701860 219085 701861
rect 219019 701796 219020 701860
rect 219084 701796 219085 701860
rect 219019 701795 219085 701796
rect 219203 701860 219269 701861
rect 219203 701796 219204 701860
rect 219268 701796 219269 701860
rect 219203 701795 219269 701796
rect 226379 701860 226445 701861
rect 226379 701796 226380 701860
rect 226444 701796 226445 701860
rect 226379 701795 226445 701796
rect 219022 700909 219082 701795
rect 219019 700908 219085 700909
rect 219019 700844 219020 700908
rect 219084 700844 219085 700908
rect 219019 700843 219085 700844
rect 215339 280804 215405 280805
rect 215339 280740 215340 280804
rect 215404 280740 215405 280804
rect 215339 280739 215405 280740
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 277174 204134 279792
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 244894 207854 279792
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 248614 211574 279792
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 255454 218414 281792
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 219206 205730 219266 701795
rect 226382 280941 226442 701795
rect 234662 700365 234722 702339
rect 235794 701792 236414 705242
rect 239514 703792 240134 707162
rect 243234 703792 243854 709082
rect 246954 703792 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 237419 702404 237485 702405
rect 237419 702340 237420 702404
rect 237484 702340 237485 702404
rect 237419 702339 237485 702340
rect 234659 700364 234725 700365
rect 234659 700300 234660 700364
rect 234724 700300 234725 700364
rect 234659 700299 234725 700300
rect 228440 687454 228760 687486
rect 228440 687218 228482 687454
rect 228718 687218 228760 687454
rect 228440 687134 228760 687218
rect 228440 686898 228482 687134
rect 228718 686898 228760 687134
rect 228440 686866 228760 686898
rect 228440 651454 228760 651486
rect 228440 651218 228482 651454
rect 228718 651218 228760 651454
rect 228440 651134 228760 651218
rect 228440 650898 228482 651134
rect 228718 650898 228760 651134
rect 228440 650866 228760 650898
rect 228440 615454 228760 615486
rect 228440 615218 228482 615454
rect 228718 615218 228760 615454
rect 228440 615134 228760 615218
rect 228440 614898 228482 615134
rect 228718 614898 228760 615134
rect 228440 614866 228760 614898
rect 228440 579454 228760 579486
rect 228440 579218 228482 579454
rect 228718 579218 228760 579454
rect 228440 579134 228760 579218
rect 228440 578898 228482 579134
rect 228718 578898 228760 579134
rect 228440 578866 228760 578898
rect 228440 543454 228760 543486
rect 228440 543218 228482 543454
rect 228718 543218 228760 543454
rect 228440 543134 228760 543218
rect 228440 542898 228482 543134
rect 228718 542898 228760 543134
rect 228440 542866 228760 542898
rect 228440 507454 228760 507486
rect 228440 507218 228482 507454
rect 228718 507218 228760 507454
rect 228440 507134 228760 507218
rect 228440 506898 228482 507134
rect 228718 506898 228760 507134
rect 228440 506866 228760 506898
rect 228440 471454 228760 471486
rect 228440 471218 228482 471454
rect 228718 471218 228760 471454
rect 228440 471134 228760 471218
rect 228440 470898 228482 471134
rect 228718 470898 228760 471134
rect 228440 470866 228760 470898
rect 228440 435454 228760 435486
rect 228440 435218 228482 435454
rect 228718 435218 228760 435454
rect 228440 435134 228760 435218
rect 228440 434898 228482 435134
rect 228718 434898 228760 435134
rect 228440 434866 228760 434898
rect 228440 399454 228760 399486
rect 228440 399218 228482 399454
rect 228718 399218 228760 399454
rect 228440 399134 228760 399218
rect 228440 398898 228482 399134
rect 228718 398898 228760 399134
rect 228440 398866 228760 398898
rect 228440 363454 228760 363486
rect 228440 363218 228482 363454
rect 228718 363218 228760 363454
rect 228440 363134 228760 363218
rect 228440 362898 228482 363134
rect 228718 362898 228760 363134
rect 228440 362866 228760 362898
rect 228440 327454 228760 327486
rect 228440 327218 228482 327454
rect 228718 327218 228760 327454
rect 228440 327134 228760 327218
rect 228440 326898 228482 327134
rect 228718 326898 228760 327134
rect 228440 326866 228760 326898
rect 228440 291454 228760 291486
rect 228440 291218 228482 291454
rect 228718 291218 228760 291454
rect 228440 291134 228760 291218
rect 228440 290898 228482 291134
rect 228718 290898 228760 291134
rect 228440 290866 228760 290898
rect 226379 280940 226445 280941
rect 226379 280876 226380 280940
rect 226444 280876 226445 280940
rect 226379 280875 226445 280876
rect 221514 259174 222134 279792
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 219387 205732 219453 205733
rect 219387 205730 219388 205732
rect 219206 205670 219388 205730
rect 219387 205668 219388 205670
rect 219452 205668 219453 205732
rect 219387 205667 219453 205668
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 262894 225854 279792
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 266614 229574 279792
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 273454 236414 281792
rect 237422 280805 237482 702339
rect 244779 702268 244845 702269
rect 244779 702204 244780 702268
rect 244844 702204 244845 702268
rect 244779 702203 244845 702204
rect 243800 669454 244120 669486
rect 243800 669218 243842 669454
rect 244078 669218 244120 669454
rect 243800 669134 244120 669218
rect 243800 668898 243842 669134
rect 244078 668898 244120 669134
rect 243800 668866 244120 668898
rect 243800 633454 244120 633486
rect 243800 633218 243842 633454
rect 244078 633218 244120 633454
rect 243800 633134 244120 633218
rect 243800 632898 243842 633134
rect 244078 632898 244120 633134
rect 243800 632866 244120 632898
rect 243800 597454 244120 597486
rect 243800 597218 243842 597454
rect 244078 597218 244120 597454
rect 243800 597134 244120 597218
rect 243800 596898 243842 597134
rect 244078 596898 244120 597134
rect 243800 596866 244120 596898
rect 243800 561454 244120 561486
rect 243800 561218 243842 561454
rect 244078 561218 244120 561454
rect 243800 561134 244120 561218
rect 243800 560898 243842 561134
rect 244078 560898 244120 561134
rect 243800 560866 244120 560898
rect 243800 525454 244120 525486
rect 243800 525218 243842 525454
rect 244078 525218 244120 525454
rect 243800 525134 244120 525218
rect 243800 524898 243842 525134
rect 244078 524898 244120 525134
rect 243800 524866 244120 524898
rect 243800 489454 244120 489486
rect 243800 489218 243842 489454
rect 244078 489218 244120 489454
rect 243800 489134 244120 489218
rect 243800 488898 243842 489134
rect 244078 488898 244120 489134
rect 243800 488866 244120 488898
rect 243800 453454 244120 453486
rect 243800 453218 243842 453454
rect 244078 453218 244120 453454
rect 243800 453134 244120 453218
rect 243800 452898 243842 453134
rect 244078 452898 244120 453134
rect 243800 452866 244120 452898
rect 243800 417454 244120 417486
rect 243800 417218 243842 417454
rect 244078 417218 244120 417454
rect 243800 417134 244120 417218
rect 243800 416898 243842 417134
rect 244078 416898 244120 417134
rect 243800 416866 244120 416898
rect 243800 381454 244120 381486
rect 243800 381218 243842 381454
rect 244078 381218 244120 381454
rect 243800 381134 244120 381218
rect 243800 380898 243842 381134
rect 244078 380898 244120 381134
rect 243800 380866 244120 380898
rect 243800 345454 244120 345486
rect 243800 345218 243842 345454
rect 244078 345218 244120 345454
rect 243800 345134 244120 345218
rect 243800 344898 243842 345134
rect 244078 344898 244120 345134
rect 243800 344866 244120 344898
rect 243800 309454 244120 309486
rect 243800 309218 243842 309454
rect 244078 309218 244120 309454
rect 243800 309134 244120 309218
rect 243800 308898 243842 309134
rect 244078 308898 244120 309134
rect 243800 308866 244120 308898
rect 237419 280804 237485 280805
rect 237419 280740 237420 280804
rect 237484 280740 237485 280804
rect 237419 280739 237485 280740
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 277174 240134 279792
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 244894 243854 279792
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 244782 191861 244842 702203
rect 247723 701996 247789 701997
rect 247723 701932 247724 701996
rect 247788 701932 247789 701996
rect 247723 701931 247789 701932
rect 246954 248614 247574 279792
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 244779 191860 244845 191861
rect 244779 191796 244780 191860
rect 244844 191796 244845 191860
rect 244779 191795 244845 191796
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 247726 165749 247786 701931
rect 253794 701792 254414 704282
rect 257514 703792 258134 706202
rect 261234 703792 261854 708122
rect 264954 703792 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 701792 272414 705242
rect 275514 703792 276134 707162
rect 279234 703792 279854 709082
rect 282954 703792 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 701792 290414 704282
rect 293514 703792 294134 706202
rect 297234 703792 297854 708122
rect 300954 703792 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 701792 308414 705242
rect 311514 703792 312134 707162
rect 315234 703792 315854 709082
rect 318954 703792 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 324267 703628 324333 703629
rect 324267 703564 324268 703628
rect 324332 703564 324333 703628
rect 324267 703563 324333 703564
rect 311755 702540 311821 702541
rect 311755 702476 311756 702540
rect 311820 702476 311821 702540
rect 311755 702475 311821 702476
rect 311758 700909 311818 702475
rect 312307 702268 312373 702269
rect 312307 702204 312308 702268
rect 312372 702204 312373 702268
rect 312307 702203 312373 702204
rect 311755 700908 311821 700909
rect 311755 700844 311756 700908
rect 311820 700844 311821 700908
rect 311755 700843 311821 700844
rect 312310 700501 312370 702203
rect 324270 701045 324330 703563
rect 325794 701792 326414 704282
rect 329514 703792 330134 706202
rect 333234 703792 333854 708122
rect 336954 703792 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 342851 702540 342917 702541
rect 342851 702476 342852 702540
rect 342916 702476 342917 702540
rect 342851 702475 342917 702476
rect 327027 702268 327093 702269
rect 327027 702204 327028 702268
rect 327092 702204 327093 702268
rect 327027 702203 327093 702204
rect 324267 701044 324333 701045
rect 324267 700980 324268 701044
rect 324332 700980 324333 701044
rect 324267 700979 324333 700980
rect 327030 700637 327090 702203
rect 342854 701045 342914 702475
rect 343794 701792 344414 705242
rect 347514 703792 348134 707162
rect 351234 703792 351854 709082
rect 354954 703792 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 354627 702540 354693 702541
rect 354627 702476 354628 702540
rect 354692 702476 354693 702540
rect 354627 702475 354693 702476
rect 355179 702540 355245 702541
rect 355179 702476 355180 702540
rect 355244 702476 355245 702540
rect 355179 702475 355245 702476
rect 360331 702540 360397 702541
rect 360331 702476 360332 702540
rect 360396 702476 360397 702540
rect 360331 702475 360397 702476
rect 354630 702130 354690 702475
rect 354630 702070 354874 702130
rect 342851 701044 342917 701045
rect 342851 700980 342852 701044
rect 342916 700980 342917 701044
rect 342851 700979 342917 700980
rect 354814 700909 354874 702070
rect 355182 701045 355242 702475
rect 357939 702132 358005 702133
rect 357939 702068 357940 702132
rect 358004 702068 358005 702132
rect 357939 702067 358005 702068
rect 360147 702132 360213 702133
rect 360147 702068 360148 702132
rect 360212 702130 360213 702132
rect 360334 702130 360394 702475
rect 360212 702070 360394 702130
rect 360212 702068 360213 702070
rect 360147 702067 360213 702068
rect 355179 701044 355245 701045
rect 355179 700980 355180 701044
rect 355244 700980 355245 701044
rect 355179 700979 355245 700980
rect 354811 700908 354877 700909
rect 354811 700844 354812 700908
rect 354876 700844 354877 700908
rect 354811 700843 354877 700844
rect 327027 700636 327093 700637
rect 327027 700572 327028 700636
rect 327092 700572 327093 700636
rect 327027 700571 327093 700572
rect 312307 700500 312373 700501
rect 312307 700436 312308 700500
rect 312372 700436 312373 700500
rect 312307 700435 312373 700436
rect 259160 687454 259480 687486
rect 259160 687218 259202 687454
rect 259438 687218 259480 687454
rect 259160 687134 259480 687218
rect 259160 686898 259202 687134
rect 259438 686898 259480 687134
rect 259160 686866 259480 686898
rect 289880 687454 290200 687486
rect 289880 687218 289922 687454
rect 290158 687218 290200 687454
rect 289880 687134 290200 687218
rect 289880 686898 289922 687134
rect 290158 686898 290200 687134
rect 289880 686866 290200 686898
rect 320600 687454 320920 687486
rect 320600 687218 320642 687454
rect 320878 687218 320920 687454
rect 320600 687134 320920 687218
rect 320600 686898 320642 687134
rect 320878 686898 320920 687134
rect 320600 686866 320920 686898
rect 351320 687454 351640 687486
rect 351320 687218 351362 687454
rect 351598 687218 351640 687454
rect 351320 687134 351640 687218
rect 351320 686898 351362 687134
rect 351598 686898 351640 687134
rect 351320 686866 351640 686898
rect 274520 669454 274840 669486
rect 274520 669218 274562 669454
rect 274798 669218 274840 669454
rect 274520 669134 274840 669218
rect 274520 668898 274562 669134
rect 274798 668898 274840 669134
rect 274520 668866 274840 668898
rect 305240 669454 305560 669486
rect 305240 669218 305282 669454
rect 305518 669218 305560 669454
rect 305240 669134 305560 669218
rect 305240 668898 305282 669134
rect 305518 668898 305560 669134
rect 305240 668866 305560 668898
rect 335960 669454 336280 669486
rect 335960 669218 336002 669454
rect 336238 669218 336280 669454
rect 335960 669134 336280 669218
rect 335960 668898 336002 669134
rect 336238 668898 336280 669134
rect 335960 668866 336280 668898
rect 259160 651454 259480 651486
rect 259160 651218 259202 651454
rect 259438 651218 259480 651454
rect 259160 651134 259480 651218
rect 259160 650898 259202 651134
rect 259438 650898 259480 651134
rect 259160 650866 259480 650898
rect 289880 651454 290200 651486
rect 289880 651218 289922 651454
rect 290158 651218 290200 651454
rect 289880 651134 290200 651218
rect 289880 650898 289922 651134
rect 290158 650898 290200 651134
rect 289880 650866 290200 650898
rect 320600 651454 320920 651486
rect 320600 651218 320642 651454
rect 320878 651218 320920 651454
rect 320600 651134 320920 651218
rect 320600 650898 320642 651134
rect 320878 650898 320920 651134
rect 320600 650866 320920 650898
rect 351320 651454 351640 651486
rect 351320 651218 351362 651454
rect 351598 651218 351640 651454
rect 351320 651134 351640 651218
rect 351320 650898 351362 651134
rect 351598 650898 351640 651134
rect 351320 650866 351640 650898
rect 274520 633454 274840 633486
rect 274520 633218 274562 633454
rect 274798 633218 274840 633454
rect 274520 633134 274840 633218
rect 274520 632898 274562 633134
rect 274798 632898 274840 633134
rect 274520 632866 274840 632898
rect 305240 633454 305560 633486
rect 305240 633218 305282 633454
rect 305518 633218 305560 633454
rect 305240 633134 305560 633218
rect 305240 632898 305282 633134
rect 305518 632898 305560 633134
rect 305240 632866 305560 632898
rect 335960 633454 336280 633486
rect 335960 633218 336002 633454
rect 336238 633218 336280 633454
rect 335960 633134 336280 633218
rect 335960 632898 336002 633134
rect 336238 632898 336280 633134
rect 335960 632866 336280 632898
rect 259160 615454 259480 615486
rect 259160 615218 259202 615454
rect 259438 615218 259480 615454
rect 259160 615134 259480 615218
rect 259160 614898 259202 615134
rect 259438 614898 259480 615134
rect 259160 614866 259480 614898
rect 289880 615454 290200 615486
rect 289880 615218 289922 615454
rect 290158 615218 290200 615454
rect 289880 615134 290200 615218
rect 289880 614898 289922 615134
rect 290158 614898 290200 615134
rect 289880 614866 290200 614898
rect 320600 615454 320920 615486
rect 320600 615218 320642 615454
rect 320878 615218 320920 615454
rect 320600 615134 320920 615218
rect 320600 614898 320642 615134
rect 320878 614898 320920 615134
rect 320600 614866 320920 614898
rect 351320 615454 351640 615486
rect 351320 615218 351362 615454
rect 351598 615218 351640 615454
rect 351320 615134 351640 615218
rect 351320 614898 351362 615134
rect 351598 614898 351640 615134
rect 351320 614866 351640 614898
rect 274520 597454 274840 597486
rect 274520 597218 274562 597454
rect 274798 597218 274840 597454
rect 274520 597134 274840 597218
rect 274520 596898 274562 597134
rect 274798 596898 274840 597134
rect 274520 596866 274840 596898
rect 305240 597454 305560 597486
rect 305240 597218 305282 597454
rect 305518 597218 305560 597454
rect 305240 597134 305560 597218
rect 305240 596898 305282 597134
rect 305518 596898 305560 597134
rect 305240 596866 305560 596898
rect 335960 597454 336280 597486
rect 335960 597218 336002 597454
rect 336238 597218 336280 597454
rect 335960 597134 336280 597218
rect 335960 596898 336002 597134
rect 336238 596898 336280 597134
rect 335960 596866 336280 596898
rect 259160 579454 259480 579486
rect 259160 579218 259202 579454
rect 259438 579218 259480 579454
rect 259160 579134 259480 579218
rect 259160 578898 259202 579134
rect 259438 578898 259480 579134
rect 259160 578866 259480 578898
rect 289880 579454 290200 579486
rect 289880 579218 289922 579454
rect 290158 579218 290200 579454
rect 289880 579134 290200 579218
rect 289880 578898 289922 579134
rect 290158 578898 290200 579134
rect 289880 578866 290200 578898
rect 320600 579454 320920 579486
rect 320600 579218 320642 579454
rect 320878 579218 320920 579454
rect 320600 579134 320920 579218
rect 320600 578898 320642 579134
rect 320878 578898 320920 579134
rect 320600 578866 320920 578898
rect 351320 579454 351640 579486
rect 351320 579218 351362 579454
rect 351598 579218 351640 579454
rect 351320 579134 351640 579218
rect 351320 578898 351362 579134
rect 351598 578898 351640 579134
rect 351320 578866 351640 578898
rect 274520 561454 274840 561486
rect 274520 561218 274562 561454
rect 274798 561218 274840 561454
rect 274520 561134 274840 561218
rect 274520 560898 274562 561134
rect 274798 560898 274840 561134
rect 274520 560866 274840 560898
rect 305240 561454 305560 561486
rect 305240 561218 305282 561454
rect 305518 561218 305560 561454
rect 305240 561134 305560 561218
rect 305240 560898 305282 561134
rect 305518 560898 305560 561134
rect 305240 560866 305560 560898
rect 335960 561454 336280 561486
rect 335960 561218 336002 561454
rect 336238 561218 336280 561454
rect 335960 561134 336280 561218
rect 335960 560898 336002 561134
rect 336238 560898 336280 561134
rect 335960 560866 336280 560898
rect 259160 543454 259480 543486
rect 259160 543218 259202 543454
rect 259438 543218 259480 543454
rect 259160 543134 259480 543218
rect 259160 542898 259202 543134
rect 259438 542898 259480 543134
rect 259160 542866 259480 542898
rect 289880 543454 290200 543486
rect 289880 543218 289922 543454
rect 290158 543218 290200 543454
rect 289880 543134 290200 543218
rect 289880 542898 289922 543134
rect 290158 542898 290200 543134
rect 289880 542866 290200 542898
rect 320600 543454 320920 543486
rect 320600 543218 320642 543454
rect 320878 543218 320920 543454
rect 320600 543134 320920 543218
rect 320600 542898 320642 543134
rect 320878 542898 320920 543134
rect 320600 542866 320920 542898
rect 351320 543454 351640 543486
rect 351320 543218 351362 543454
rect 351598 543218 351640 543454
rect 351320 543134 351640 543218
rect 351320 542898 351362 543134
rect 351598 542898 351640 543134
rect 351320 542866 351640 542898
rect 274520 525454 274840 525486
rect 274520 525218 274562 525454
rect 274798 525218 274840 525454
rect 274520 525134 274840 525218
rect 274520 524898 274562 525134
rect 274798 524898 274840 525134
rect 274520 524866 274840 524898
rect 305240 525454 305560 525486
rect 305240 525218 305282 525454
rect 305518 525218 305560 525454
rect 305240 525134 305560 525218
rect 305240 524898 305282 525134
rect 305518 524898 305560 525134
rect 305240 524866 305560 524898
rect 335960 525454 336280 525486
rect 335960 525218 336002 525454
rect 336238 525218 336280 525454
rect 335960 525134 336280 525218
rect 335960 524898 336002 525134
rect 336238 524898 336280 525134
rect 335960 524866 336280 524898
rect 259160 507454 259480 507486
rect 259160 507218 259202 507454
rect 259438 507218 259480 507454
rect 259160 507134 259480 507218
rect 259160 506898 259202 507134
rect 259438 506898 259480 507134
rect 259160 506866 259480 506898
rect 289880 507454 290200 507486
rect 289880 507218 289922 507454
rect 290158 507218 290200 507454
rect 289880 507134 290200 507218
rect 289880 506898 289922 507134
rect 290158 506898 290200 507134
rect 289880 506866 290200 506898
rect 320600 507454 320920 507486
rect 320600 507218 320642 507454
rect 320878 507218 320920 507454
rect 320600 507134 320920 507218
rect 320600 506898 320642 507134
rect 320878 506898 320920 507134
rect 320600 506866 320920 506898
rect 351320 507454 351640 507486
rect 351320 507218 351362 507454
rect 351598 507218 351640 507454
rect 351320 507134 351640 507218
rect 351320 506898 351362 507134
rect 351598 506898 351640 507134
rect 351320 506866 351640 506898
rect 274520 489454 274840 489486
rect 274520 489218 274562 489454
rect 274798 489218 274840 489454
rect 274520 489134 274840 489218
rect 274520 488898 274562 489134
rect 274798 488898 274840 489134
rect 274520 488866 274840 488898
rect 305240 489454 305560 489486
rect 305240 489218 305282 489454
rect 305518 489218 305560 489454
rect 305240 489134 305560 489218
rect 305240 488898 305282 489134
rect 305518 488898 305560 489134
rect 305240 488866 305560 488898
rect 335960 489454 336280 489486
rect 335960 489218 336002 489454
rect 336238 489218 336280 489454
rect 335960 489134 336280 489218
rect 335960 488898 336002 489134
rect 336238 488898 336280 489134
rect 335960 488866 336280 488898
rect 259160 471454 259480 471486
rect 259160 471218 259202 471454
rect 259438 471218 259480 471454
rect 259160 471134 259480 471218
rect 259160 470898 259202 471134
rect 259438 470898 259480 471134
rect 259160 470866 259480 470898
rect 289880 471454 290200 471486
rect 289880 471218 289922 471454
rect 290158 471218 290200 471454
rect 289880 471134 290200 471218
rect 289880 470898 289922 471134
rect 290158 470898 290200 471134
rect 289880 470866 290200 470898
rect 320600 471454 320920 471486
rect 320600 471218 320642 471454
rect 320878 471218 320920 471454
rect 320600 471134 320920 471218
rect 320600 470898 320642 471134
rect 320878 470898 320920 471134
rect 320600 470866 320920 470898
rect 351320 471454 351640 471486
rect 351320 471218 351362 471454
rect 351598 471218 351640 471454
rect 351320 471134 351640 471218
rect 351320 470898 351362 471134
rect 351598 470898 351640 471134
rect 351320 470866 351640 470898
rect 274520 453454 274840 453486
rect 274520 453218 274562 453454
rect 274798 453218 274840 453454
rect 274520 453134 274840 453218
rect 274520 452898 274562 453134
rect 274798 452898 274840 453134
rect 274520 452866 274840 452898
rect 305240 453454 305560 453486
rect 305240 453218 305282 453454
rect 305518 453218 305560 453454
rect 305240 453134 305560 453218
rect 305240 452898 305282 453134
rect 305518 452898 305560 453134
rect 305240 452866 305560 452898
rect 335960 453454 336280 453486
rect 335960 453218 336002 453454
rect 336238 453218 336280 453454
rect 335960 453134 336280 453218
rect 335960 452898 336002 453134
rect 336238 452898 336280 453134
rect 335960 452866 336280 452898
rect 259160 435454 259480 435486
rect 259160 435218 259202 435454
rect 259438 435218 259480 435454
rect 259160 435134 259480 435218
rect 259160 434898 259202 435134
rect 259438 434898 259480 435134
rect 259160 434866 259480 434898
rect 289880 435454 290200 435486
rect 289880 435218 289922 435454
rect 290158 435218 290200 435454
rect 289880 435134 290200 435218
rect 289880 434898 289922 435134
rect 290158 434898 290200 435134
rect 289880 434866 290200 434898
rect 320600 435454 320920 435486
rect 320600 435218 320642 435454
rect 320878 435218 320920 435454
rect 320600 435134 320920 435218
rect 320600 434898 320642 435134
rect 320878 434898 320920 435134
rect 320600 434866 320920 434898
rect 351320 435454 351640 435486
rect 351320 435218 351362 435454
rect 351598 435218 351640 435454
rect 351320 435134 351640 435218
rect 351320 434898 351362 435134
rect 351598 434898 351640 435134
rect 351320 434866 351640 434898
rect 274520 417454 274840 417486
rect 274520 417218 274562 417454
rect 274798 417218 274840 417454
rect 274520 417134 274840 417218
rect 274520 416898 274562 417134
rect 274798 416898 274840 417134
rect 274520 416866 274840 416898
rect 305240 417454 305560 417486
rect 305240 417218 305282 417454
rect 305518 417218 305560 417454
rect 305240 417134 305560 417218
rect 305240 416898 305282 417134
rect 305518 416898 305560 417134
rect 305240 416866 305560 416898
rect 335960 417454 336280 417486
rect 335960 417218 336002 417454
rect 336238 417218 336280 417454
rect 335960 417134 336280 417218
rect 335960 416898 336002 417134
rect 336238 416898 336280 417134
rect 335960 416866 336280 416898
rect 259160 399454 259480 399486
rect 259160 399218 259202 399454
rect 259438 399218 259480 399454
rect 259160 399134 259480 399218
rect 259160 398898 259202 399134
rect 259438 398898 259480 399134
rect 259160 398866 259480 398898
rect 289880 399454 290200 399486
rect 289880 399218 289922 399454
rect 290158 399218 290200 399454
rect 289880 399134 290200 399218
rect 289880 398898 289922 399134
rect 290158 398898 290200 399134
rect 289880 398866 290200 398898
rect 320600 399454 320920 399486
rect 320600 399218 320642 399454
rect 320878 399218 320920 399454
rect 320600 399134 320920 399218
rect 320600 398898 320642 399134
rect 320878 398898 320920 399134
rect 320600 398866 320920 398898
rect 351320 399454 351640 399486
rect 351320 399218 351362 399454
rect 351598 399218 351640 399454
rect 351320 399134 351640 399218
rect 351320 398898 351362 399134
rect 351598 398898 351640 399134
rect 351320 398866 351640 398898
rect 274520 381454 274840 381486
rect 274520 381218 274562 381454
rect 274798 381218 274840 381454
rect 274520 381134 274840 381218
rect 274520 380898 274562 381134
rect 274798 380898 274840 381134
rect 274520 380866 274840 380898
rect 305240 381454 305560 381486
rect 305240 381218 305282 381454
rect 305518 381218 305560 381454
rect 305240 381134 305560 381218
rect 305240 380898 305282 381134
rect 305518 380898 305560 381134
rect 305240 380866 305560 380898
rect 335960 381454 336280 381486
rect 335960 381218 336002 381454
rect 336238 381218 336280 381454
rect 335960 381134 336280 381218
rect 335960 380898 336002 381134
rect 336238 380898 336280 381134
rect 335960 380866 336280 380898
rect 259160 363454 259480 363486
rect 259160 363218 259202 363454
rect 259438 363218 259480 363454
rect 259160 363134 259480 363218
rect 259160 362898 259202 363134
rect 259438 362898 259480 363134
rect 259160 362866 259480 362898
rect 289880 363454 290200 363486
rect 289880 363218 289922 363454
rect 290158 363218 290200 363454
rect 289880 363134 290200 363218
rect 289880 362898 289922 363134
rect 290158 362898 290200 363134
rect 289880 362866 290200 362898
rect 320600 363454 320920 363486
rect 320600 363218 320642 363454
rect 320878 363218 320920 363454
rect 320600 363134 320920 363218
rect 320600 362898 320642 363134
rect 320878 362898 320920 363134
rect 320600 362866 320920 362898
rect 351320 363454 351640 363486
rect 351320 363218 351362 363454
rect 351598 363218 351640 363454
rect 351320 363134 351640 363218
rect 351320 362898 351362 363134
rect 351598 362898 351640 363134
rect 351320 362866 351640 362898
rect 274520 345454 274840 345486
rect 274520 345218 274562 345454
rect 274798 345218 274840 345454
rect 274520 345134 274840 345218
rect 274520 344898 274562 345134
rect 274798 344898 274840 345134
rect 274520 344866 274840 344898
rect 305240 345454 305560 345486
rect 305240 345218 305282 345454
rect 305518 345218 305560 345454
rect 305240 345134 305560 345218
rect 305240 344898 305282 345134
rect 305518 344898 305560 345134
rect 305240 344866 305560 344898
rect 335960 345454 336280 345486
rect 335960 345218 336002 345454
rect 336238 345218 336280 345454
rect 335960 345134 336280 345218
rect 335960 344898 336002 345134
rect 336238 344898 336280 345134
rect 335960 344866 336280 344898
rect 259160 327454 259480 327486
rect 259160 327218 259202 327454
rect 259438 327218 259480 327454
rect 259160 327134 259480 327218
rect 259160 326898 259202 327134
rect 259438 326898 259480 327134
rect 259160 326866 259480 326898
rect 289880 327454 290200 327486
rect 289880 327218 289922 327454
rect 290158 327218 290200 327454
rect 289880 327134 290200 327218
rect 289880 326898 289922 327134
rect 290158 326898 290200 327134
rect 289880 326866 290200 326898
rect 320600 327454 320920 327486
rect 320600 327218 320642 327454
rect 320878 327218 320920 327454
rect 320600 327134 320920 327218
rect 320600 326898 320642 327134
rect 320878 326898 320920 327134
rect 320600 326866 320920 326898
rect 351320 327454 351640 327486
rect 351320 327218 351362 327454
rect 351598 327218 351640 327454
rect 351320 327134 351640 327218
rect 351320 326898 351362 327134
rect 351598 326898 351640 327134
rect 351320 326866 351640 326898
rect 274520 309454 274840 309486
rect 274520 309218 274562 309454
rect 274798 309218 274840 309454
rect 274520 309134 274840 309218
rect 274520 308898 274562 309134
rect 274798 308898 274840 309134
rect 274520 308866 274840 308898
rect 305240 309454 305560 309486
rect 305240 309218 305282 309454
rect 305518 309218 305560 309454
rect 305240 309134 305560 309218
rect 305240 308898 305282 309134
rect 305518 308898 305560 309134
rect 305240 308866 305560 308898
rect 335960 309454 336280 309486
rect 335960 309218 336002 309454
rect 336238 309218 336280 309454
rect 335960 309134 336280 309218
rect 335960 308898 336002 309134
rect 336238 308898 336280 309134
rect 335960 308866 336280 308898
rect 259160 291454 259480 291486
rect 259160 291218 259202 291454
rect 259438 291218 259480 291454
rect 259160 291134 259480 291218
rect 259160 290898 259202 291134
rect 259438 290898 259480 291134
rect 259160 290866 259480 290898
rect 289880 291454 290200 291486
rect 289880 291218 289922 291454
rect 290158 291218 290200 291454
rect 289880 291134 290200 291218
rect 289880 290898 289922 291134
rect 290158 290898 290200 291134
rect 289880 290866 290200 290898
rect 320600 291454 320920 291486
rect 320600 291218 320642 291454
rect 320878 291218 320920 291454
rect 320600 291134 320920 291218
rect 320600 290898 320642 291134
rect 320878 290898 320920 291134
rect 320600 290866 320920 290898
rect 351320 291454 351640 291486
rect 351320 291218 351362 291454
rect 351598 291218 351640 291454
rect 351320 291134 351640 291218
rect 351320 290898 351362 291134
rect 351598 290898 351640 291134
rect 351320 290866 351640 290898
rect 253794 255454 254414 281792
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 247723 165748 247789 165749
rect 247723 165684 247724 165748
rect 247788 165684 247789 165748
rect 247723 165683 247789 165684
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 259174 258134 279792
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 262894 261854 279792
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 266614 265574 279792
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 273454 272414 281792
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 277174 276134 279792
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 244894 279854 279792
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 248614 283574 279792
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 255454 290414 281792
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 259174 294134 279792
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 262894 297854 279792
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 266614 301574 279792
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 273454 308414 281792
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 277174 312134 279792
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 244894 315854 279792
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 248614 319574 279792
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 255454 326414 281792
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 259174 330134 279792
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 262894 333854 279792
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 266614 337574 279792
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 273454 344414 281792
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 277174 348134 279792
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 244894 351854 279792
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 248614 355574 279792
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 357942 99517 358002 702067
rect 361794 701792 362414 704282
rect 365514 703792 366134 706202
rect 366955 703900 367021 703901
rect 366955 703836 366956 703900
rect 367020 703836 367021 703900
rect 366955 703835 367021 703836
rect 365667 702540 365733 702541
rect 365667 702476 365668 702540
rect 365732 702476 365733 702540
rect 365667 702475 365733 702476
rect 365670 700773 365730 702475
rect 366958 701450 367018 703835
rect 369234 703792 369854 708122
rect 372954 703792 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 701792 380414 705242
rect 383514 703792 384134 707162
rect 387234 703792 387854 709082
rect 390954 703792 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 701792 398414 704282
rect 401514 703792 402134 706202
rect 405234 703792 405854 708122
rect 408954 703792 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 701792 416414 705242
rect 419514 703792 420134 707162
rect 423234 703792 423854 709082
rect 426954 703792 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 419395 702540 419461 702541
rect 419395 702476 419396 702540
rect 419460 702476 419461 702540
rect 419395 702475 419461 702476
rect 366958 701390 367570 701450
rect 367510 701045 367570 701390
rect 367507 701044 367573 701045
rect 367507 700980 367508 701044
rect 367572 700980 367573 701044
rect 367507 700979 367573 700980
rect 419398 700773 419458 702475
rect 433794 701792 434414 704282
rect 437514 703792 438134 706202
rect 441234 703792 441854 708122
rect 444954 703792 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 701792 452414 705242
rect 455514 703792 456134 707162
rect 459234 703792 459854 709082
rect 462954 703792 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 701792 470414 704282
rect 473514 703792 474134 706202
rect 477234 703792 477854 708122
rect 480954 703792 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 481035 702540 481101 702541
rect 481035 702476 481036 702540
rect 481100 702476 481101 702540
rect 481035 702475 481101 702476
rect 365667 700772 365733 700773
rect 365667 700708 365668 700772
rect 365732 700708 365733 700772
rect 365667 700707 365733 700708
rect 419395 700772 419461 700773
rect 419395 700708 419396 700772
rect 419460 700708 419461 700772
rect 419395 700707 419461 700708
rect 481038 700093 481098 702475
rect 487794 701792 488414 705242
rect 491514 703792 492134 707162
rect 495234 703792 495854 709082
rect 498954 703792 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 701792 506414 704282
rect 509514 703792 510134 706202
rect 513234 703792 513854 708122
rect 516954 703792 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 701792 524414 705242
rect 527514 703792 528134 707162
rect 531234 703792 531854 709082
rect 534954 703792 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 701792 542414 704282
rect 545514 703792 546134 706202
rect 549234 703792 549854 708122
rect 552954 703792 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 701792 560414 705242
rect 563514 703792 564134 707162
rect 567234 703792 567854 709082
rect 570954 703792 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577267 703220 577333 703221
rect 577267 703156 577268 703220
rect 577332 703156 577333 703220
rect 577267 703155 577333 703156
rect 577083 702540 577149 702541
rect 577083 702476 577084 702540
rect 577148 702476 577149 702540
rect 577083 702475 577149 702476
rect 574691 702404 574757 702405
rect 574691 702340 574692 702404
rect 574756 702340 574757 702404
rect 574691 702339 574757 702340
rect 494651 701316 494717 701317
rect 494651 701252 494652 701316
rect 494716 701252 494717 701316
rect 494651 701251 494717 701252
rect 506427 701316 506493 701317
rect 506427 701252 506428 701316
rect 506492 701252 506493 701316
rect 506427 701251 506493 701252
rect 494654 700909 494714 701251
rect 494651 700908 494717 700909
rect 494651 700844 494652 700908
rect 494716 700844 494717 700908
rect 494651 700843 494717 700844
rect 481035 700092 481101 700093
rect 481035 700028 481036 700092
rect 481100 700028 481101 700092
rect 481035 700027 481101 700028
rect 382040 687454 382360 687486
rect 382040 687218 382082 687454
rect 382318 687218 382360 687454
rect 382040 687134 382360 687218
rect 382040 686898 382082 687134
rect 382318 686898 382360 687134
rect 382040 686866 382360 686898
rect 412760 687454 413080 687486
rect 412760 687218 412802 687454
rect 413038 687218 413080 687454
rect 412760 687134 413080 687218
rect 412760 686898 412802 687134
rect 413038 686898 413080 687134
rect 412760 686866 413080 686898
rect 443480 687454 443800 687486
rect 443480 687218 443522 687454
rect 443758 687218 443800 687454
rect 443480 687134 443800 687218
rect 443480 686898 443522 687134
rect 443758 686898 443800 687134
rect 443480 686866 443800 686898
rect 474200 687454 474520 687486
rect 474200 687218 474242 687454
rect 474478 687218 474520 687454
rect 474200 687134 474520 687218
rect 474200 686898 474242 687134
rect 474478 686898 474520 687134
rect 474200 686866 474520 686898
rect 504920 687454 505240 687486
rect 504920 687218 504962 687454
rect 505198 687218 505240 687454
rect 504920 687134 505240 687218
rect 504920 686898 504962 687134
rect 505198 686898 505240 687134
rect 504920 686866 505240 686898
rect 366680 669454 367000 669486
rect 366680 669218 366722 669454
rect 366958 669218 367000 669454
rect 366680 669134 367000 669218
rect 366680 668898 366722 669134
rect 366958 668898 367000 669134
rect 366680 668866 367000 668898
rect 397400 669454 397720 669486
rect 397400 669218 397442 669454
rect 397678 669218 397720 669454
rect 397400 669134 397720 669218
rect 397400 668898 397442 669134
rect 397678 668898 397720 669134
rect 397400 668866 397720 668898
rect 428120 669454 428440 669486
rect 428120 669218 428162 669454
rect 428398 669218 428440 669454
rect 428120 669134 428440 669218
rect 428120 668898 428162 669134
rect 428398 668898 428440 669134
rect 428120 668866 428440 668898
rect 458840 669454 459160 669486
rect 458840 669218 458882 669454
rect 459118 669218 459160 669454
rect 458840 669134 459160 669218
rect 458840 668898 458882 669134
rect 459118 668898 459160 669134
rect 458840 668866 459160 668898
rect 489560 669454 489880 669486
rect 489560 669218 489602 669454
rect 489838 669218 489880 669454
rect 489560 669134 489880 669218
rect 489560 668898 489602 669134
rect 489838 668898 489880 669134
rect 489560 668866 489880 668898
rect 382040 651454 382360 651486
rect 382040 651218 382082 651454
rect 382318 651218 382360 651454
rect 382040 651134 382360 651218
rect 382040 650898 382082 651134
rect 382318 650898 382360 651134
rect 382040 650866 382360 650898
rect 412760 651454 413080 651486
rect 412760 651218 412802 651454
rect 413038 651218 413080 651454
rect 412760 651134 413080 651218
rect 412760 650898 412802 651134
rect 413038 650898 413080 651134
rect 412760 650866 413080 650898
rect 443480 651454 443800 651486
rect 443480 651218 443522 651454
rect 443758 651218 443800 651454
rect 443480 651134 443800 651218
rect 443480 650898 443522 651134
rect 443758 650898 443800 651134
rect 443480 650866 443800 650898
rect 474200 651454 474520 651486
rect 474200 651218 474242 651454
rect 474478 651218 474520 651454
rect 474200 651134 474520 651218
rect 474200 650898 474242 651134
rect 474478 650898 474520 651134
rect 474200 650866 474520 650898
rect 504920 651454 505240 651486
rect 504920 651218 504962 651454
rect 505198 651218 505240 651454
rect 504920 651134 505240 651218
rect 504920 650898 504962 651134
rect 505198 650898 505240 651134
rect 504920 650866 505240 650898
rect 366680 633454 367000 633486
rect 366680 633218 366722 633454
rect 366958 633218 367000 633454
rect 366680 633134 367000 633218
rect 366680 632898 366722 633134
rect 366958 632898 367000 633134
rect 366680 632866 367000 632898
rect 397400 633454 397720 633486
rect 397400 633218 397442 633454
rect 397678 633218 397720 633454
rect 397400 633134 397720 633218
rect 397400 632898 397442 633134
rect 397678 632898 397720 633134
rect 397400 632866 397720 632898
rect 428120 633454 428440 633486
rect 428120 633218 428162 633454
rect 428398 633218 428440 633454
rect 428120 633134 428440 633218
rect 428120 632898 428162 633134
rect 428398 632898 428440 633134
rect 428120 632866 428440 632898
rect 458840 633454 459160 633486
rect 458840 633218 458882 633454
rect 459118 633218 459160 633454
rect 458840 633134 459160 633218
rect 458840 632898 458882 633134
rect 459118 632898 459160 633134
rect 458840 632866 459160 632898
rect 489560 633454 489880 633486
rect 489560 633218 489602 633454
rect 489838 633218 489880 633454
rect 489560 633134 489880 633218
rect 489560 632898 489602 633134
rect 489838 632898 489880 633134
rect 489560 632866 489880 632898
rect 382040 615454 382360 615486
rect 382040 615218 382082 615454
rect 382318 615218 382360 615454
rect 382040 615134 382360 615218
rect 382040 614898 382082 615134
rect 382318 614898 382360 615134
rect 382040 614866 382360 614898
rect 412760 615454 413080 615486
rect 412760 615218 412802 615454
rect 413038 615218 413080 615454
rect 412760 615134 413080 615218
rect 412760 614898 412802 615134
rect 413038 614898 413080 615134
rect 412760 614866 413080 614898
rect 443480 615454 443800 615486
rect 443480 615218 443522 615454
rect 443758 615218 443800 615454
rect 443480 615134 443800 615218
rect 443480 614898 443522 615134
rect 443758 614898 443800 615134
rect 443480 614866 443800 614898
rect 474200 615454 474520 615486
rect 474200 615218 474242 615454
rect 474478 615218 474520 615454
rect 474200 615134 474520 615218
rect 474200 614898 474242 615134
rect 474478 614898 474520 615134
rect 474200 614866 474520 614898
rect 504920 615454 505240 615486
rect 504920 615218 504962 615454
rect 505198 615218 505240 615454
rect 504920 615134 505240 615218
rect 504920 614898 504962 615134
rect 505198 614898 505240 615134
rect 504920 614866 505240 614898
rect 366680 597454 367000 597486
rect 366680 597218 366722 597454
rect 366958 597218 367000 597454
rect 366680 597134 367000 597218
rect 366680 596898 366722 597134
rect 366958 596898 367000 597134
rect 366680 596866 367000 596898
rect 397400 597454 397720 597486
rect 397400 597218 397442 597454
rect 397678 597218 397720 597454
rect 397400 597134 397720 597218
rect 397400 596898 397442 597134
rect 397678 596898 397720 597134
rect 397400 596866 397720 596898
rect 428120 597454 428440 597486
rect 428120 597218 428162 597454
rect 428398 597218 428440 597454
rect 428120 597134 428440 597218
rect 428120 596898 428162 597134
rect 428398 596898 428440 597134
rect 428120 596866 428440 596898
rect 458840 597454 459160 597486
rect 458840 597218 458882 597454
rect 459118 597218 459160 597454
rect 458840 597134 459160 597218
rect 458840 596898 458882 597134
rect 459118 596898 459160 597134
rect 458840 596866 459160 596898
rect 489560 597454 489880 597486
rect 489560 597218 489602 597454
rect 489838 597218 489880 597454
rect 489560 597134 489880 597218
rect 489560 596898 489602 597134
rect 489838 596898 489880 597134
rect 489560 596866 489880 596898
rect 382040 579454 382360 579486
rect 382040 579218 382082 579454
rect 382318 579218 382360 579454
rect 382040 579134 382360 579218
rect 382040 578898 382082 579134
rect 382318 578898 382360 579134
rect 382040 578866 382360 578898
rect 412760 579454 413080 579486
rect 412760 579218 412802 579454
rect 413038 579218 413080 579454
rect 412760 579134 413080 579218
rect 412760 578898 412802 579134
rect 413038 578898 413080 579134
rect 412760 578866 413080 578898
rect 443480 579454 443800 579486
rect 443480 579218 443522 579454
rect 443758 579218 443800 579454
rect 443480 579134 443800 579218
rect 443480 578898 443522 579134
rect 443758 578898 443800 579134
rect 443480 578866 443800 578898
rect 474200 579454 474520 579486
rect 474200 579218 474242 579454
rect 474478 579218 474520 579454
rect 474200 579134 474520 579218
rect 474200 578898 474242 579134
rect 474478 578898 474520 579134
rect 474200 578866 474520 578898
rect 504920 579454 505240 579486
rect 504920 579218 504962 579454
rect 505198 579218 505240 579454
rect 504920 579134 505240 579218
rect 504920 578898 504962 579134
rect 505198 578898 505240 579134
rect 504920 578866 505240 578898
rect 366680 561454 367000 561486
rect 366680 561218 366722 561454
rect 366958 561218 367000 561454
rect 366680 561134 367000 561218
rect 366680 560898 366722 561134
rect 366958 560898 367000 561134
rect 366680 560866 367000 560898
rect 397400 561454 397720 561486
rect 397400 561218 397442 561454
rect 397678 561218 397720 561454
rect 397400 561134 397720 561218
rect 397400 560898 397442 561134
rect 397678 560898 397720 561134
rect 397400 560866 397720 560898
rect 428120 561454 428440 561486
rect 428120 561218 428162 561454
rect 428398 561218 428440 561454
rect 428120 561134 428440 561218
rect 428120 560898 428162 561134
rect 428398 560898 428440 561134
rect 428120 560866 428440 560898
rect 458840 561454 459160 561486
rect 458840 561218 458882 561454
rect 459118 561218 459160 561454
rect 458840 561134 459160 561218
rect 458840 560898 458882 561134
rect 459118 560898 459160 561134
rect 458840 560866 459160 560898
rect 489560 561454 489880 561486
rect 489560 561218 489602 561454
rect 489838 561218 489880 561454
rect 489560 561134 489880 561218
rect 489560 560898 489602 561134
rect 489838 560898 489880 561134
rect 489560 560866 489880 560898
rect 382040 543454 382360 543486
rect 382040 543218 382082 543454
rect 382318 543218 382360 543454
rect 382040 543134 382360 543218
rect 382040 542898 382082 543134
rect 382318 542898 382360 543134
rect 382040 542866 382360 542898
rect 412760 543454 413080 543486
rect 412760 543218 412802 543454
rect 413038 543218 413080 543454
rect 412760 543134 413080 543218
rect 412760 542898 412802 543134
rect 413038 542898 413080 543134
rect 412760 542866 413080 542898
rect 443480 543454 443800 543486
rect 443480 543218 443522 543454
rect 443758 543218 443800 543454
rect 443480 543134 443800 543218
rect 443480 542898 443522 543134
rect 443758 542898 443800 543134
rect 443480 542866 443800 542898
rect 474200 543454 474520 543486
rect 474200 543218 474242 543454
rect 474478 543218 474520 543454
rect 474200 543134 474520 543218
rect 474200 542898 474242 543134
rect 474478 542898 474520 543134
rect 474200 542866 474520 542898
rect 504920 543454 505240 543486
rect 504920 543218 504962 543454
rect 505198 543218 505240 543454
rect 504920 543134 505240 543218
rect 504920 542898 504962 543134
rect 505198 542898 505240 543134
rect 504920 542866 505240 542898
rect 366680 525454 367000 525486
rect 366680 525218 366722 525454
rect 366958 525218 367000 525454
rect 366680 525134 367000 525218
rect 366680 524898 366722 525134
rect 366958 524898 367000 525134
rect 366680 524866 367000 524898
rect 397400 525454 397720 525486
rect 397400 525218 397442 525454
rect 397678 525218 397720 525454
rect 397400 525134 397720 525218
rect 397400 524898 397442 525134
rect 397678 524898 397720 525134
rect 397400 524866 397720 524898
rect 428120 525454 428440 525486
rect 428120 525218 428162 525454
rect 428398 525218 428440 525454
rect 428120 525134 428440 525218
rect 428120 524898 428162 525134
rect 428398 524898 428440 525134
rect 428120 524866 428440 524898
rect 458840 525454 459160 525486
rect 458840 525218 458882 525454
rect 459118 525218 459160 525454
rect 458840 525134 459160 525218
rect 458840 524898 458882 525134
rect 459118 524898 459160 525134
rect 458840 524866 459160 524898
rect 489560 525454 489880 525486
rect 489560 525218 489602 525454
rect 489838 525218 489880 525454
rect 489560 525134 489880 525218
rect 489560 524898 489602 525134
rect 489838 524898 489880 525134
rect 489560 524866 489880 524898
rect 382040 507454 382360 507486
rect 382040 507218 382082 507454
rect 382318 507218 382360 507454
rect 382040 507134 382360 507218
rect 382040 506898 382082 507134
rect 382318 506898 382360 507134
rect 382040 506866 382360 506898
rect 412760 507454 413080 507486
rect 412760 507218 412802 507454
rect 413038 507218 413080 507454
rect 412760 507134 413080 507218
rect 412760 506898 412802 507134
rect 413038 506898 413080 507134
rect 412760 506866 413080 506898
rect 443480 507454 443800 507486
rect 443480 507218 443522 507454
rect 443758 507218 443800 507454
rect 443480 507134 443800 507218
rect 443480 506898 443522 507134
rect 443758 506898 443800 507134
rect 443480 506866 443800 506898
rect 474200 507454 474520 507486
rect 474200 507218 474242 507454
rect 474478 507218 474520 507454
rect 474200 507134 474520 507218
rect 474200 506898 474242 507134
rect 474478 506898 474520 507134
rect 474200 506866 474520 506898
rect 504920 507454 505240 507486
rect 504920 507218 504962 507454
rect 505198 507218 505240 507454
rect 504920 507134 505240 507218
rect 504920 506898 504962 507134
rect 505198 506898 505240 507134
rect 504920 506866 505240 506898
rect 366680 489454 367000 489486
rect 366680 489218 366722 489454
rect 366958 489218 367000 489454
rect 366680 489134 367000 489218
rect 366680 488898 366722 489134
rect 366958 488898 367000 489134
rect 366680 488866 367000 488898
rect 397400 489454 397720 489486
rect 397400 489218 397442 489454
rect 397678 489218 397720 489454
rect 397400 489134 397720 489218
rect 397400 488898 397442 489134
rect 397678 488898 397720 489134
rect 397400 488866 397720 488898
rect 428120 489454 428440 489486
rect 428120 489218 428162 489454
rect 428398 489218 428440 489454
rect 428120 489134 428440 489218
rect 428120 488898 428162 489134
rect 428398 488898 428440 489134
rect 428120 488866 428440 488898
rect 458840 489454 459160 489486
rect 458840 489218 458882 489454
rect 459118 489218 459160 489454
rect 458840 489134 459160 489218
rect 458840 488898 458882 489134
rect 459118 488898 459160 489134
rect 458840 488866 459160 488898
rect 489560 489454 489880 489486
rect 489560 489218 489602 489454
rect 489838 489218 489880 489454
rect 489560 489134 489880 489218
rect 489560 488898 489602 489134
rect 489838 488898 489880 489134
rect 489560 488866 489880 488898
rect 382040 471454 382360 471486
rect 382040 471218 382082 471454
rect 382318 471218 382360 471454
rect 382040 471134 382360 471218
rect 382040 470898 382082 471134
rect 382318 470898 382360 471134
rect 382040 470866 382360 470898
rect 412760 471454 413080 471486
rect 412760 471218 412802 471454
rect 413038 471218 413080 471454
rect 412760 471134 413080 471218
rect 412760 470898 412802 471134
rect 413038 470898 413080 471134
rect 412760 470866 413080 470898
rect 443480 471454 443800 471486
rect 443480 471218 443522 471454
rect 443758 471218 443800 471454
rect 443480 471134 443800 471218
rect 443480 470898 443522 471134
rect 443758 470898 443800 471134
rect 443480 470866 443800 470898
rect 474200 471454 474520 471486
rect 474200 471218 474242 471454
rect 474478 471218 474520 471454
rect 474200 471134 474520 471218
rect 474200 470898 474242 471134
rect 474478 470898 474520 471134
rect 474200 470866 474520 470898
rect 504920 471454 505240 471486
rect 504920 471218 504962 471454
rect 505198 471218 505240 471454
rect 504920 471134 505240 471218
rect 504920 470898 504962 471134
rect 505198 470898 505240 471134
rect 504920 470866 505240 470898
rect 366680 453454 367000 453486
rect 366680 453218 366722 453454
rect 366958 453218 367000 453454
rect 366680 453134 367000 453218
rect 366680 452898 366722 453134
rect 366958 452898 367000 453134
rect 366680 452866 367000 452898
rect 397400 453454 397720 453486
rect 397400 453218 397442 453454
rect 397678 453218 397720 453454
rect 397400 453134 397720 453218
rect 397400 452898 397442 453134
rect 397678 452898 397720 453134
rect 397400 452866 397720 452898
rect 428120 453454 428440 453486
rect 428120 453218 428162 453454
rect 428398 453218 428440 453454
rect 428120 453134 428440 453218
rect 428120 452898 428162 453134
rect 428398 452898 428440 453134
rect 428120 452866 428440 452898
rect 458840 453454 459160 453486
rect 458840 453218 458882 453454
rect 459118 453218 459160 453454
rect 458840 453134 459160 453218
rect 458840 452898 458882 453134
rect 459118 452898 459160 453134
rect 458840 452866 459160 452898
rect 489560 453454 489880 453486
rect 489560 453218 489602 453454
rect 489838 453218 489880 453454
rect 489560 453134 489880 453218
rect 489560 452898 489602 453134
rect 489838 452898 489880 453134
rect 489560 452866 489880 452898
rect 382040 435454 382360 435486
rect 382040 435218 382082 435454
rect 382318 435218 382360 435454
rect 382040 435134 382360 435218
rect 382040 434898 382082 435134
rect 382318 434898 382360 435134
rect 382040 434866 382360 434898
rect 412760 435454 413080 435486
rect 412760 435218 412802 435454
rect 413038 435218 413080 435454
rect 412760 435134 413080 435218
rect 412760 434898 412802 435134
rect 413038 434898 413080 435134
rect 412760 434866 413080 434898
rect 443480 435454 443800 435486
rect 443480 435218 443522 435454
rect 443758 435218 443800 435454
rect 443480 435134 443800 435218
rect 443480 434898 443522 435134
rect 443758 434898 443800 435134
rect 443480 434866 443800 434898
rect 474200 435454 474520 435486
rect 474200 435218 474242 435454
rect 474478 435218 474520 435454
rect 474200 435134 474520 435218
rect 474200 434898 474242 435134
rect 474478 434898 474520 435134
rect 474200 434866 474520 434898
rect 504920 435454 505240 435486
rect 504920 435218 504962 435454
rect 505198 435218 505240 435454
rect 504920 435134 505240 435218
rect 504920 434898 504962 435134
rect 505198 434898 505240 435134
rect 504920 434866 505240 434898
rect 366680 417454 367000 417486
rect 366680 417218 366722 417454
rect 366958 417218 367000 417454
rect 366680 417134 367000 417218
rect 366680 416898 366722 417134
rect 366958 416898 367000 417134
rect 366680 416866 367000 416898
rect 397400 417454 397720 417486
rect 397400 417218 397442 417454
rect 397678 417218 397720 417454
rect 397400 417134 397720 417218
rect 397400 416898 397442 417134
rect 397678 416898 397720 417134
rect 397400 416866 397720 416898
rect 428120 417454 428440 417486
rect 428120 417218 428162 417454
rect 428398 417218 428440 417454
rect 428120 417134 428440 417218
rect 428120 416898 428162 417134
rect 428398 416898 428440 417134
rect 428120 416866 428440 416898
rect 458840 417454 459160 417486
rect 458840 417218 458882 417454
rect 459118 417218 459160 417454
rect 458840 417134 459160 417218
rect 458840 416898 458882 417134
rect 459118 416898 459160 417134
rect 458840 416866 459160 416898
rect 489560 417454 489880 417486
rect 489560 417218 489602 417454
rect 489838 417218 489880 417454
rect 489560 417134 489880 417218
rect 489560 416898 489602 417134
rect 489838 416898 489880 417134
rect 489560 416866 489880 416898
rect 382040 399454 382360 399486
rect 382040 399218 382082 399454
rect 382318 399218 382360 399454
rect 382040 399134 382360 399218
rect 382040 398898 382082 399134
rect 382318 398898 382360 399134
rect 382040 398866 382360 398898
rect 412760 399454 413080 399486
rect 412760 399218 412802 399454
rect 413038 399218 413080 399454
rect 412760 399134 413080 399218
rect 412760 398898 412802 399134
rect 413038 398898 413080 399134
rect 412760 398866 413080 398898
rect 443480 399454 443800 399486
rect 443480 399218 443522 399454
rect 443758 399218 443800 399454
rect 443480 399134 443800 399218
rect 443480 398898 443522 399134
rect 443758 398898 443800 399134
rect 443480 398866 443800 398898
rect 474200 399454 474520 399486
rect 474200 399218 474242 399454
rect 474478 399218 474520 399454
rect 474200 399134 474520 399218
rect 474200 398898 474242 399134
rect 474478 398898 474520 399134
rect 474200 398866 474520 398898
rect 504920 399454 505240 399486
rect 504920 399218 504962 399454
rect 505198 399218 505240 399454
rect 504920 399134 505240 399218
rect 504920 398898 504962 399134
rect 505198 398898 505240 399134
rect 504920 398866 505240 398898
rect 366680 381454 367000 381486
rect 366680 381218 366722 381454
rect 366958 381218 367000 381454
rect 366680 381134 367000 381218
rect 366680 380898 366722 381134
rect 366958 380898 367000 381134
rect 366680 380866 367000 380898
rect 397400 381454 397720 381486
rect 397400 381218 397442 381454
rect 397678 381218 397720 381454
rect 397400 381134 397720 381218
rect 397400 380898 397442 381134
rect 397678 380898 397720 381134
rect 397400 380866 397720 380898
rect 428120 381454 428440 381486
rect 428120 381218 428162 381454
rect 428398 381218 428440 381454
rect 428120 381134 428440 381218
rect 428120 380898 428162 381134
rect 428398 380898 428440 381134
rect 428120 380866 428440 380898
rect 458840 381454 459160 381486
rect 458840 381218 458882 381454
rect 459118 381218 459160 381454
rect 458840 381134 459160 381218
rect 458840 380898 458882 381134
rect 459118 380898 459160 381134
rect 458840 380866 459160 380898
rect 489560 381454 489880 381486
rect 489560 381218 489602 381454
rect 489838 381218 489880 381454
rect 489560 381134 489880 381218
rect 489560 380898 489602 381134
rect 489838 380898 489880 381134
rect 489560 380866 489880 380898
rect 382040 363454 382360 363486
rect 382040 363218 382082 363454
rect 382318 363218 382360 363454
rect 382040 363134 382360 363218
rect 382040 362898 382082 363134
rect 382318 362898 382360 363134
rect 382040 362866 382360 362898
rect 412760 363454 413080 363486
rect 412760 363218 412802 363454
rect 413038 363218 413080 363454
rect 412760 363134 413080 363218
rect 412760 362898 412802 363134
rect 413038 362898 413080 363134
rect 412760 362866 413080 362898
rect 443480 363454 443800 363486
rect 443480 363218 443522 363454
rect 443758 363218 443800 363454
rect 443480 363134 443800 363218
rect 443480 362898 443522 363134
rect 443758 362898 443800 363134
rect 443480 362866 443800 362898
rect 474200 363454 474520 363486
rect 474200 363218 474242 363454
rect 474478 363218 474520 363454
rect 474200 363134 474520 363218
rect 474200 362898 474242 363134
rect 474478 362898 474520 363134
rect 474200 362866 474520 362898
rect 504920 363454 505240 363486
rect 504920 363218 504962 363454
rect 505198 363218 505240 363454
rect 504920 363134 505240 363218
rect 504920 362898 504962 363134
rect 505198 362898 505240 363134
rect 504920 362866 505240 362898
rect 366680 345454 367000 345486
rect 366680 345218 366722 345454
rect 366958 345218 367000 345454
rect 366680 345134 367000 345218
rect 366680 344898 366722 345134
rect 366958 344898 367000 345134
rect 366680 344866 367000 344898
rect 397400 345454 397720 345486
rect 397400 345218 397442 345454
rect 397678 345218 397720 345454
rect 397400 345134 397720 345218
rect 397400 344898 397442 345134
rect 397678 344898 397720 345134
rect 397400 344866 397720 344898
rect 428120 345454 428440 345486
rect 428120 345218 428162 345454
rect 428398 345218 428440 345454
rect 428120 345134 428440 345218
rect 428120 344898 428162 345134
rect 428398 344898 428440 345134
rect 428120 344866 428440 344898
rect 458840 345454 459160 345486
rect 458840 345218 458882 345454
rect 459118 345218 459160 345454
rect 458840 345134 459160 345218
rect 458840 344898 458882 345134
rect 459118 344898 459160 345134
rect 458840 344866 459160 344898
rect 489560 345454 489880 345486
rect 489560 345218 489602 345454
rect 489838 345218 489880 345454
rect 489560 345134 489880 345218
rect 489560 344898 489602 345134
rect 489838 344898 489880 345134
rect 489560 344866 489880 344898
rect 382040 327454 382360 327486
rect 382040 327218 382082 327454
rect 382318 327218 382360 327454
rect 382040 327134 382360 327218
rect 382040 326898 382082 327134
rect 382318 326898 382360 327134
rect 382040 326866 382360 326898
rect 412760 327454 413080 327486
rect 412760 327218 412802 327454
rect 413038 327218 413080 327454
rect 412760 327134 413080 327218
rect 412760 326898 412802 327134
rect 413038 326898 413080 327134
rect 412760 326866 413080 326898
rect 443480 327454 443800 327486
rect 443480 327218 443522 327454
rect 443758 327218 443800 327454
rect 443480 327134 443800 327218
rect 443480 326898 443522 327134
rect 443758 326898 443800 327134
rect 443480 326866 443800 326898
rect 474200 327454 474520 327486
rect 474200 327218 474242 327454
rect 474478 327218 474520 327454
rect 474200 327134 474520 327218
rect 474200 326898 474242 327134
rect 474478 326898 474520 327134
rect 474200 326866 474520 326898
rect 504920 327454 505240 327486
rect 504920 327218 504962 327454
rect 505198 327218 505240 327454
rect 504920 327134 505240 327218
rect 504920 326898 504962 327134
rect 505198 326898 505240 327134
rect 504920 326866 505240 326898
rect 366680 309454 367000 309486
rect 366680 309218 366722 309454
rect 366958 309218 367000 309454
rect 366680 309134 367000 309218
rect 366680 308898 366722 309134
rect 366958 308898 367000 309134
rect 366680 308866 367000 308898
rect 397400 309454 397720 309486
rect 397400 309218 397442 309454
rect 397678 309218 397720 309454
rect 397400 309134 397720 309218
rect 397400 308898 397442 309134
rect 397678 308898 397720 309134
rect 397400 308866 397720 308898
rect 428120 309454 428440 309486
rect 428120 309218 428162 309454
rect 428398 309218 428440 309454
rect 428120 309134 428440 309218
rect 428120 308898 428162 309134
rect 428398 308898 428440 309134
rect 428120 308866 428440 308898
rect 458840 309454 459160 309486
rect 458840 309218 458882 309454
rect 459118 309218 459160 309454
rect 458840 309134 459160 309218
rect 458840 308898 458882 309134
rect 459118 308898 459160 309134
rect 458840 308866 459160 308898
rect 489560 309454 489880 309486
rect 489560 309218 489602 309454
rect 489838 309218 489880 309454
rect 489560 309134 489880 309218
rect 489560 308898 489602 309134
rect 489838 308898 489880 309134
rect 489560 308866 489880 308898
rect 382040 291454 382360 291486
rect 382040 291218 382082 291454
rect 382318 291218 382360 291454
rect 382040 291134 382360 291218
rect 382040 290898 382082 291134
rect 382318 290898 382360 291134
rect 382040 290866 382360 290898
rect 412760 291454 413080 291486
rect 412760 291218 412802 291454
rect 413038 291218 413080 291454
rect 412760 291134 413080 291218
rect 412760 290898 412802 291134
rect 413038 290898 413080 291134
rect 412760 290866 413080 290898
rect 443480 291454 443800 291486
rect 443480 291218 443522 291454
rect 443758 291218 443800 291454
rect 443480 291134 443800 291218
rect 443480 290898 443522 291134
rect 443758 290898 443800 291134
rect 443480 290866 443800 290898
rect 474200 291454 474520 291486
rect 474200 291218 474242 291454
rect 474478 291218 474520 291454
rect 474200 291134 474520 291218
rect 474200 290898 474242 291134
rect 474478 290898 474520 291134
rect 474200 290866 474520 290898
rect 504920 291454 505240 291486
rect 504920 291218 504962 291454
rect 505198 291218 505240 291454
rect 504920 291134 505240 291218
rect 504920 290898 504962 291134
rect 505198 290898 505240 291134
rect 504920 290866 505240 290898
rect 506430 283797 506490 701251
rect 517651 701180 517717 701181
rect 517651 701116 517652 701180
rect 517716 701116 517717 701180
rect 517651 701115 517717 701116
rect 521699 701180 521765 701181
rect 521699 701116 521700 701180
rect 521764 701116 521765 701180
rect 521699 701115 521765 701116
rect 525379 701180 525445 701181
rect 525379 701116 525380 701180
rect 525444 701116 525445 701180
rect 525379 701115 525445 701116
rect 528323 701180 528389 701181
rect 528323 701116 528324 701180
rect 528388 701116 528389 701180
rect 528323 701115 528389 701116
rect 533291 701180 533357 701181
rect 533291 701116 533292 701180
rect 533356 701116 533357 701180
rect 533291 701115 533357 701116
rect 572667 701180 572733 701181
rect 572667 701116 572668 701180
rect 572732 701116 572733 701180
rect 572667 701115 572733 701116
rect 517654 287070 517714 701115
rect 521702 699821 521762 701115
rect 525382 699957 525442 701115
rect 525379 699956 525445 699957
rect 525379 699892 525380 699956
rect 525444 699892 525445 699956
rect 525379 699891 525445 699892
rect 521699 699820 521765 699821
rect 521699 699756 521700 699820
rect 521764 699756 521765 699820
rect 521699 699755 521765 699756
rect 520280 669454 520600 669486
rect 520280 669218 520322 669454
rect 520558 669218 520600 669454
rect 520280 669134 520600 669218
rect 520280 668898 520322 669134
rect 520558 668898 520600 669134
rect 520280 668866 520600 668898
rect 520280 633454 520600 633486
rect 520280 633218 520322 633454
rect 520558 633218 520600 633454
rect 520280 633134 520600 633218
rect 520280 632898 520322 633134
rect 520558 632898 520600 633134
rect 520280 632866 520600 632898
rect 520280 597454 520600 597486
rect 520280 597218 520322 597454
rect 520558 597218 520600 597454
rect 520280 597134 520600 597218
rect 520280 596898 520322 597134
rect 520558 596898 520600 597134
rect 520280 596866 520600 596898
rect 520280 561454 520600 561486
rect 520280 561218 520322 561454
rect 520558 561218 520600 561454
rect 520280 561134 520600 561218
rect 520280 560898 520322 561134
rect 520558 560898 520600 561134
rect 520280 560866 520600 560898
rect 520280 525454 520600 525486
rect 520280 525218 520322 525454
rect 520558 525218 520600 525454
rect 520280 525134 520600 525218
rect 520280 524898 520322 525134
rect 520558 524898 520600 525134
rect 520280 524866 520600 524898
rect 520280 489454 520600 489486
rect 520280 489218 520322 489454
rect 520558 489218 520600 489454
rect 520280 489134 520600 489218
rect 520280 488898 520322 489134
rect 520558 488898 520600 489134
rect 520280 488866 520600 488898
rect 520280 453454 520600 453486
rect 520280 453218 520322 453454
rect 520558 453218 520600 453454
rect 520280 453134 520600 453218
rect 520280 452898 520322 453134
rect 520558 452898 520600 453134
rect 520280 452866 520600 452898
rect 520280 417454 520600 417486
rect 520280 417218 520322 417454
rect 520558 417218 520600 417454
rect 520280 417134 520600 417218
rect 520280 416898 520322 417134
rect 520558 416898 520600 417134
rect 520280 416866 520600 416898
rect 520280 381454 520600 381486
rect 520280 381218 520322 381454
rect 520558 381218 520600 381454
rect 520280 381134 520600 381218
rect 520280 380898 520322 381134
rect 520558 380898 520600 381134
rect 520280 380866 520600 380898
rect 520280 345454 520600 345486
rect 520280 345218 520322 345454
rect 520558 345218 520600 345454
rect 520280 345134 520600 345218
rect 520280 344898 520322 345134
rect 520558 344898 520600 345134
rect 520280 344866 520600 344898
rect 520280 309454 520600 309486
rect 520280 309218 520322 309454
rect 520558 309218 520600 309454
rect 520280 309134 520600 309218
rect 520280 308898 520322 309134
rect 520558 308898 520600 309134
rect 520280 308866 520600 308898
rect 517654 287010 517898 287070
rect 506427 283796 506493 283797
rect 506427 283732 506428 283796
rect 506492 283732 506493 283796
rect 506427 283731 506493 283732
rect 361794 255454 362414 281792
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 357939 99516 358005 99517
rect 357939 99452 357940 99516
rect 358004 99452 358005 99516
rect 357939 99451 358005 99452
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 259174 366134 279792
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 262894 369854 279792
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 266614 373574 279792
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 273454 380414 281792
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 277174 384134 279792
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 244894 387854 279792
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 248614 391574 279792
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 255454 398414 281792
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 259174 402134 279792
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 262894 405854 279792
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 266614 409574 279792
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 273454 416414 281792
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 277174 420134 279792
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 244894 423854 279792
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 248614 427574 279792
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 255454 434414 281792
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 259174 438134 279792
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 262894 441854 279792
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 266614 445574 279792
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 273454 452414 281792
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 277174 456134 279792
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 244894 459854 279792
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 248614 463574 279792
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 255454 470414 281792
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 259174 474134 279792
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 262894 477854 279792
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 266614 481574 279792
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 273454 488414 281792
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 277174 492134 279792
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 244894 495854 279792
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 248614 499574 279792
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 255454 506414 281792
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 259174 510134 279792
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 262894 513854 279792
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 266614 517574 279792
rect 517838 267749 517898 287010
rect 523794 273454 524414 281792
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 517835 267748 517901 267749
rect 517835 267684 517836 267748
rect 517900 267684 517901 267748
rect 517835 267683 517901 267684
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 277174 528134 279792
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 528326 215253 528386 701115
rect 531234 244894 531854 279792
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 528323 215252 528389 215253
rect 528323 215188 528324 215252
rect 528388 215188 528389 215252
rect 528323 215187 528389 215188
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 533294 202877 533354 701115
rect 535640 687454 535960 687486
rect 535640 687218 535682 687454
rect 535918 687218 535960 687454
rect 535640 687134 535960 687218
rect 535640 686898 535682 687134
rect 535918 686898 535960 687134
rect 535640 686866 535960 686898
rect 566360 687454 566680 687486
rect 566360 687218 566402 687454
rect 566638 687218 566680 687454
rect 566360 687134 566680 687218
rect 566360 686898 566402 687134
rect 566638 686898 566680 687134
rect 566360 686866 566680 686898
rect 551000 669454 551320 669486
rect 551000 669218 551042 669454
rect 551278 669218 551320 669454
rect 551000 669134 551320 669218
rect 551000 668898 551042 669134
rect 551278 668898 551320 669134
rect 551000 668866 551320 668898
rect 535640 651454 535960 651486
rect 535640 651218 535682 651454
rect 535918 651218 535960 651454
rect 535640 651134 535960 651218
rect 535640 650898 535682 651134
rect 535918 650898 535960 651134
rect 535640 650866 535960 650898
rect 566360 651454 566680 651486
rect 566360 651218 566402 651454
rect 566638 651218 566680 651454
rect 566360 651134 566680 651218
rect 566360 650898 566402 651134
rect 566638 650898 566680 651134
rect 566360 650866 566680 650898
rect 551000 633454 551320 633486
rect 551000 633218 551042 633454
rect 551278 633218 551320 633454
rect 551000 633134 551320 633218
rect 551000 632898 551042 633134
rect 551278 632898 551320 633134
rect 551000 632866 551320 632898
rect 535640 615454 535960 615486
rect 535640 615218 535682 615454
rect 535918 615218 535960 615454
rect 535640 615134 535960 615218
rect 535640 614898 535682 615134
rect 535918 614898 535960 615134
rect 535640 614866 535960 614898
rect 566360 615454 566680 615486
rect 566360 615218 566402 615454
rect 566638 615218 566680 615454
rect 566360 615134 566680 615218
rect 566360 614898 566402 615134
rect 566638 614898 566680 615134
rect 566360 614866 566680 614898
rect 551000 597454 551320 597486
rect 551000 597218 551042 597454
rect 551278 597218 551320 597454
rect 551000 597134 551320 597218
rect 551000 596898 551042 597134
rect 551278 596898 551320 597134
rect 551000 596866 551320 596898
rect 535640 579454 535960 579486
rect 535640 579218 535682 579454
rect 535918 579218 535960 579454
rect 535640 579134 535960 579218
rect 535640 578898 535682 579134
rect 535918 578898 535960 579134
rect 535640 578866 535960 578898
rect 566360 579454 566680 579486
rect 566360 579218 566402 579454
rect 566638 579218 566680 579454
rect 566360 579134 566680 579218
rect 566360 578898 566402 579134
rect 566638 578898 566680 579134
rect 566360 578866 566680 578898
rect 551000 561454 551320 561486
rect 551000 561218 551042 561454
rect 551278 561218 551320 561454
rect 551000 561134 551320 561218
rect 551000 560898 551042 561134
rect 551278 560898 551320 561134
rect 551000 560866 551320 560898
rect 535640 543454 535960 543486
rect 535640 543218 535682 543454
rect 535918 543218 535960 543454
rect 535640 543134 535960 543218
rect 535640 542898 535682 543134
rect 535918 542898 535960 543134
rect 535640 542866 535960 542898
rect 566360 543454 566680 543486
rect 566360 543218 566402 543454
rect 566638 543218 566680 543454
rect 566360 543134 566680 543218
rect 566360 542898 566402 543134
rect 566638 542898 566680 543134
rect 566360 542866 566680 542898
rect 551000 525454 551320 525486
rect 551000 525218 551042 525454
rect 551278 525218 551320 525454
rect 551000 525134 551320 525218
rect 551000 524898 551042 525134
rect 551278 524898 551320 525134
rect 551000 524866 551320 524898
rect 535640 507454 535960 507486
rect 535640 507218 535682 507454
rect 535918 507218 535960 507454
rect 535640 507134 535960 507218
rect 535640 506898 535682 507134
rect 535918 506898 535960 507134
rect 535640 506866 535960 506898
rect 566360 507454 566680 507486
rect 566360 507218 566402 507454
rect 566638 507218 566680 507454
rect 566360 507134 566680 507218
rect 566360 506898 566402 507134
rect 566638 506898 566680 507134
rect 566360 506866 566680 506898
rect 551000 489454 551320 489486
rect 551000 489218 551042 489454
rect 551278 489218 551320 489454
rect 551000 489134 551320 489218
rect 551000 488898 551042 489134
rect 551278 488898 551320 489134
rect 551000 488866 551320 488898
rect 535640 471454 535960 471486
rect 535640 471218 535682 471454
rect 535918 471218 535960 471454
rect 535640 471134 535960 471218
rect 535640 470898 535682 471134
rect 535918 470898 535960 471134
rect 535640 470866 535960 470898
rect 566360 471454 566680 471486
rect 566360 471218 566402 471454
rect 566638 471218 566680 471454
rect 566360 471134 566680 471218
rect 566360 470898 566402 471134
rect 566638 470898 566680 471134
rect 566360 470866 566680 470898
rect 551000 453454 551320 453486
rect 551000 453218 551042 453454
rect 551278 453218 551320 453454
rect 551000 453134 551320 453218
rect 551000 452898 551042 453134
rect 551278 452898 551320 453134
rect 551000 452866 551320 452898
rect 535640 435454 535960 435486
rect 535640 435218 535682 435454
rect 535918 435218 535960 435454
rect 535640 435134 535960 435218
rect 535640 434898 535682 435134
rect 535918 434898 535960 435134
rect 535640 434866 535960 434898
rect 566360 435454 566680 435486
rect 566360 435218 566402 435454
rect 566638 435218 566680 435454
rect 566360 435134 566680 435218
rect 566360 434898 566402 435134
rect 566638 434898 566680 435134
rect 566360 434866 566680 434898
rect 551000 417454 551320 417486
rect 551000 417218 551042 417454
rect 551278 417218 551320 417454
rect 551000 417134 551320 417218
rect 551000 416898 551042 417134
rect 551278 416898 551320 417134
rect 551000 416866 551320 416898
rect 535640 399454 535960 399486
rect 535640 399218 535682 399454
rect 535918 399218 535960 399454
rect 535640 399134 535960 399218
rect 535640 398898 535682 399134
rect 535918 398898 535960 399134
rect 535640 398866 535960 398898
rect 566360 399454 566680 399486
rect 566360 399218 566402 399454
rect 566638 399218 566680 399454
rect 566360 399134 566680 399218
rect 566360 398898 566402 399134
rect 566638 398898 566680 399134
rect 566360 398866 566680 398898
rect 551000 381454 551320 381486
rect 551000 381218 551042 381454
rect 551278 381218 551320 381454
rect 551000 381134 551320 381218
rect 551000 380898 551042 381134
rect 551278 380898 551320 381134
rect 551000 380866 551320 380898
rect 535640 363454 535960 363486
rect 535640 363218 535682 363454
rect 535918 363218 535960 363454
rect 535640 363134 535960 363218
rect 535640 362898 535682 363134
rect 535918 362898 535960 363134
rect 535640 362866 535960 362898
rect 566360 363454 566680 363486
rect 566360 363218 566402 363454
rect 566638 363218 566680 363454
rect 566360 363134 566680 363218
rect 566360 362898 566402 363134
rect 566638 362898 566680 363134
rect 566360 362866 566680 362898
rect 551000 345454 551320 345486
rect 551000 345218 551042 345454
rect 551278 345218 551320 345454
rect 551000 345134 551320 345218
rect 551000 344898 551042 345134
rect 551278 344898 551320 345134
rect 551000 344866 551320 344898
rect 535640 327454 535960 327486
rect 535640 327218 535682 327454
rect 535918 327218 535960 327454
rect 535640 327134 535960 327218
rect 535640 326898 535682 327134
rect 535918 326898 535960 327134
rect 535640 326866 535960 326898
rect 566360 327454 566680 327486
rect 566360 327218 566402 327454
rect 566638 327218 566680 327454
rect 566360 327134 566680 327218
rect 566360 326898 566402 327134
rect 566638 326898 566680 327134
rect 566360 326866 566680 326898
rect 551000 309454 551320 309486
rect 551000 309218 551042 309454
rect 551278 309218 551320 309454
rect 551000 309134 551320 309218
rect 551000 308898 551042 309134
rect 551278 308898 551320 309134
rect 551000 308866 551320 308898
rect 535640 291454 535960 291486
rect 535640 291218 535682 291454
rect 535918 291218 535960 291454
rect 535640 291134 535960 291218
rect 535640 290898 535682 291134
rect 535918 290898 535960 291134
rect 535640 290866 535960 290898
rect 566360 291454 566680 291486
rect 566360 291218 566402 291454
rect 566638 291218 566680 291454
rect 566360 291134 566680 291218
rect 566360 290898 566402 291134
rect 566638 290898 566680 291134
rect 566360 290866 566680 290898
rect 534954 248614 535574 279792
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 533291 202876 533357 202877
rect 533291 202812 533292 202876
rect 533356 202812 533357 202876
rect 533291 202811 533357 202812
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 255454 542414 281792
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 259174 546134 279792
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 262894 549854 279792
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 266614 553574 279792
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 273454 560414 281792
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 277174 564134 279792
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 244894 567854 279792
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 248614 571574 279792
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 572670 33149 572730 701115
rect 574694 404429 574754 702339
rect 575979 701996 576045 701997
rect 575979 701932 575980 701996
rect 576044 701932 576045 701996
rect 575979 701931 576045 701932
rect 574875 700500 574941 700501
rect 574875 700436 574876 700500
rect 574940 700436 574941 700500
rect 574875 700435 574941 700436
rect 574878 643245 574938 700435
rect 574875 643244 574941 643245
rect 574875 643180 574876 643244
rect 574940 643180 574941 643244
rect 574875 643179 574941 643180
rect 575982 591021 576042 701931
rect 575979 591020 576045 591021
rect 575979 590956 575980 591020
rect 576044 590956 576045 591020
rect 575979 590955 576045 590956
rect 577086 471477 577146 702475
rect 577083 471476 577149 471477
rect 577083 471412 577084 471476
rect 577148 471412 577149 471476
rect 577083 471411 577149 471412
rect 574691 404428 574757 404429
rect 574691 404364 574692 404428
rect 574756 404364 574757 404428
rect 574691 404363 574757 404364
rect 577270 351933 577330 703155
rect 577635 703084 577701 703085
rect 577635 703020 577636 703084
rect 577700 703020 577701 703084
rect 577635 703019 577701 703020
rect 577451 701180 577517 701181
rect 577451 701116 577452 701180
rect 577516 701116 577517 701180
rect 577451 701115 577517 701116
rect 577267 351932 577333 351933
rect 577267 351868 577268 351932
rect 577332 351868 577333 351932
rect 577267 351867 577333 351868
rect 572667 33148 572733 33149
rect 572667 33084 572668 33148
rect 572732 33084 572733 33148
rect 572667 33083 572733 33084
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577454 20637 577514 701115
rect 577638 630869 577698 703019
rect 577794 701792 578414 704282
rect 581514 703792 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 580211 703492 580277 703493
rect 580211 703428 580212 703492
rect 580276 703428 580277 703492
rect 580211 703427 580277 703428
rect 580027 703356 580093 703357
rect 580027 703292 580028 703356
rect 580092 703292 580093 703356
rect 580027 703291 580093 703292
rect 579843 700772 579909 700773
rect 579843 700708 579844 700772
rect 579908 700708 579909 700772
rect 579843 700707 579909 700708
rect 578739 700636 578805 700637
rect 578739 700572 578740 700636
rect 578804 700572 578805 700636
rect 578739 700571 578805 700572
rect 578742 683909 578802 700571
rect 579846 697237 579906 700707
rect 579843 697236 579909 697237
rect 579843 697172 579844 697236
rect 579908 697172 579909 697236
rect 579843 697171 579909 697172
rect 578739 683908 578805 683909
rect 578739 683844 578740 683908
rect 578804 683844 578805 683908
rect 578739 683843 578805 683844
rect 580030 670717 580090 703291
rect 580027 670716 580093 670717
rect 580027 670652 580028 670716
rect 580092 670652 580093 670716
rect 580027 670651 580093 670652
rect 577635 630868 577701 630869
rect 577635 630804 577636 630868
rect 577700 630804 577701 630868
rect 577635 630803 577701 630804
rect 580214 458149 580274 703427
rect 580763 702948 580829 702949
rect 580763 702884 580764 702948
rect 580828 702884 580829 702948
rect 580763 702883 580829 702884
rect 580579 702812 580645 702813
rect 580579 702748 580580 702812
rect 580644 702748 580645 702812
rect 580579 702747 580645 702748
rect 580395 702676 580461 702677
rect 580395 702612 580396 702676
rect 580460 702612 580461 702676
rect 580395 702611 580461 702612
rect 580398 511325 580458 702611
rect 580582 564365 580642 702747
rect 580766 617541 580826 702883
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 580763 617540 580829 617541
rect 580763 617476 580764 617540
rect 580828 617476 580829 617540
rect 580763 617475 580829 617476
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 580579 564364 580645 564365
rect 580579 564300 580580 564364
rect 580644 564300 580645 564364
rect 580579 564299 580645 564300
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 580395 511324 580461 511325
rect 580395 511260 580396 511324
rect 580460 511260 580461 511324
rect 580395 511259 580461 511260
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 580211 458148 580277 458149
rect 580211 458084 580212 458148
rect 580276 458084 580277 458148
rect 580211 458083 580277 458084
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 577794 255454 578414 281792
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577451 20636 577517 20637
rect 577451 20572 577452 20636
rect 577516 20572 577517 20636
rect 577451 20571 577517 20572
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 259174 582134 279792
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 167042 687218 167278 687454
rect 167042 686898 167278 687134
rect 197762 687218 197998 687454
rect 197762 686898 197998 687134
rect 182402 669218 182638 669454
rect 182402 668898 182638 669134
rect 213122 669218 213358 669454
rect 213122 668898 213358 669134
rect 167042 651218 167278 651454
rect 167042 650898 167278 651134
rect 197762 651218 197998 651454
rect 197762 650898 197998 651134
rect 182402 633218 182638 633454
rect 182402 632898 182638 633134
rect 213122 633218 213358 633454
rect 213122 632898 213358 633134
rect 167042 615218 167278 615454
rect 167042 614898 167278 615134
rect 197762 615218 197998 615454
rect 197762 614898 197998 615134
rect 182402 597218 182638 597454
rect 182402 596898 182638 597134
rect 213122 597218 213358 597454
rect 213122 596898 213358 597134
rect 167042 579218 167278 579454
rect 167042 578898 167278 579134
rect 197762 579218 197998 579454
rect 197762 578898 197998 579134
rect 182402 561218 182638 561454
rect 182402 560898 182638 561134
rect 213122 561218 213358 561454
rect 213122 560898 213358 561134
rect 167042 543218 167278 543454
rect 167042 542898 167278 543134
rect 197762 543218 197998 543454
rect 197762 542898 197998 543134
rect 182402 525218 182638 525454
rect 182402 524898 182638 525134
rect 213122 525218 213358 525454
rect 213122 524898 213358 525134
rect 167042 507218 167278 507454
rect 167042 506898 167278 507134
rect 197762 507218 197998 507454
rect 197762 506898 197998 507134
rect 182402 489218 182638 489454
rect 182402 488898 182638 489134
rect 213122 489218 213358 489454
rect 213122 488898 213358 489134
rect 167042 471218 167278 471454
rect 167042 470898 167278 471134
rect 197762 471218 197998 471454
rect 197762 470898 197998 471134
rect 182402 453218 182638 453454
rect 182402 452898 182638 453134
rect 213122 453218 213358 453454
rect 213122 452898 213358 453134
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 167042 435218 167278 435454
rect 167042 434898 167278 435134
rect 197762 435218 197998 435454
rect 197762 434898 197998 435134
rect 182402 417218 182638 417454
rect 182402 416898 182638 417134
rect 213122 417218 213358 417454
rect 213122 416898 213358 417134
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 167042 399218 167278 399454
rect 167042 398898 167278 399134
rect 197762 399218 197998 399454
rect 197762 398898 197998 399134
rect 182402 381218 182638 381454
rect 182402 380898 182638 381134
rect 213122 381218 213358 381454
rect 213122 380898 213358 381134
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 167042 363218 167278 363454
rect 167042 362898 167278 363134
rect 197762 363218 197998 363454
rect 197762 362898 197998 363134
rect 182402 345218 182638 345454
rect 182402 344898 182638 345134
rect 213122 345218 213358 345454
rect 213122 344898 213358 345134
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 167042 327218 167278 327454
rect 167042 326898 167278 327134
rect 197762 327218 197998 327454
rect 197762 326898 197998 327134
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 182402 309218 182638 309454
rect 182402 308898 182638 309134
rect 213122 309218 213358 309454
rect 213122 308898 213358 309134
rect 167042 291218 167278 291454
rect 167042 290898 167278 291134
rect 197762 291218 197998 291454
rect 197762 290898 197998 291134
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 228482 687218 228718 687454
rect 228482 686898 228718 687134
rect 228482 651218 228718 651454
rect 228482 650898 228718 651134
rect 228482 615218 228718 615454
rect 228482 614898 228718 615134
rect 228482 579218 228718 579454
rect 228482 578898 228718 579134
rect 228482 543218 228718 543454
rect 228482 542898 228718 543134
rect 228482 507218 228718 507454
rect 228482 506898 228718 507134
rect 228482 471218 228718 471454
rect 228482 470898 228718 471134
rect 228482 435218 228718 435454
rect 228482 434898 228718 435134
rect 228482 399218 228718 399454
rect 228482 398898 228718 399134
rect 228482 363218 228718 363454
rect 228482 362898 228718 363134
rect 228482 327218 228718 327454
rect 228482 326898 228718 327134
rect 228482 291218 228718 291454
rect 228482 290898 228718 291134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 243842 669218 244078 669454
rect 243842 668898 244078 669134
rect 243842 633218 244078 633454
rect 243842 632898 244078 633134
rect 243842 597218 244078 597454
rect 243842 596898 244078 597134
rect 243842 561218 244078 561454
rect 243842 560898 244078 561134
rect 243842 525218 244078 525454
rect 243842 524898 244078 525134
rect 243842 489218 244078 489454
rect 243842 488898 244078 489134
rect 243842 453218 244078 453454
rect 243842 452898 244078 453134
rect 243842 417218 244078 417454
rect 243842 416898 244078 417134
rect 243842 381218 244078 381454
rect 243842 380898 244078 381134
rect 243842 345218 244078 345454
rect 243842 344898 244078 345134
rect 243842 309218 244078 309454
rect 243842 308898 244078 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 259202 687218 259438 687454
rect 259202 686898 259438 687134
rect 289922 687218 290158 687454
rect 289922 686898 290158 687134
rect 320642 687218 320878 687454
rect 320642 686898 320878 687134
rect 351362 687218 351598 687454
rect 351362 686898 351598 687134
rect 274562 669218 274798 669454
rect 274562 668898 274798 669134
rect 305282 669218 305518 669454
rect 305282 668898 305518 669134
rect 336002 669218 336238 669454
rect 336002 668898 336238 669134
rect 259202 651218 259438 651454
rect 259202 650898 259438 651134
rect 289922 651218 290158 651454
rect 289922 650898 290158 651134
rect 320642 651218 320878 651454
rect 320642 650898 320878 651134
rect 351362 651218 351598 651454
rect 351362 650898 351598 651134
rect 274562 633218 274798 633454
rect 274562 632898 274798 633134
rect 305282 633218 305518 633454
rect 305282 632898 305518 633134
rect 336002 633218 336238 633454
rect 336002 632898 336238 633134
rect 259202 615218 259438 615454
rect 259202 614898 259438 615134
rect 289922 615218 290158 615454
rect 289922 614898 290158 615134
rect 320642 615218 320878 615454
rect 320642 614898 320878 615134
rect 351362 615218 351598 615454
rect 351362 614898 351598 615134
rect 274562 597218 274798 597454
rect 274562 596898 274798 597134
rect 305282 597218 305518 597454
rect 305282 596898 305518 597134
rect 336002 597218 336238 597454
rect 336002 596898 336238 597134
rect 259202 579218 259438 579454
rect 259202 578898 259438 579134
rect 289922 579218 290158 579454
rect 289922 578898 290158 579134
rect 320642 579218 320878 579454
rect 320642 578898 320878 579134
rect 351362 579218 351598 579454
rect 351362 578898 351598 579134
rect 274562 561218 274798 561454
rect 274562 560898 274798 561134
rect 305282 561218 305518 561454
rect 305282 560898 305518 561134
rect 336002 561218 336238 561454
rect 336002 560898 336238 561134
rect 259202 543218 259438 543454
rect 259202 542898 259438 543134
rect 289922 543218 290158 543454
rect 289922 542898 290158 543134
rect 320642 543218 320878 543454
rect 320642 542898 320878 543134
rect 351362 543218 351598 543454
rect 351362 542898 351598 543134
rect 274562 525218 274798 525454
rect 274562 524898 274798 525134
rect 305282 525218 305518 525454
rect 305282 524898 305518 525134
rect 336002 525218 336238 525454
rect 336002 524898 336238 525134
rect 259202 507218 259438 507454
rect 259202 506898 259438 507134
rect 289922 507218 290158 507454
rect 289922 506898 290158 507134
rect 320642 507218 320878 507454
rect 320642 506898 320878 507134
rect 351362 507218 351598 507454
rect 351362 506898 351598 507134
rect 274562 489218 274798 489454
rect 274562 488898 274798 489134
rect 305282 489218 305518 489454
rect 305282 488898 305518 489134
rect 336002 489218 336238 489454
rect 336002 488898 336238 489134
rect 259202 471218 259438 471454
rect 259202 470898 259438 471134
rect 289922 471218 290158 471454
rect 289922 470898 290158 471134
rect 320642 471218 320878 471454
rect 320642 470898 320878 471134
rect 351362 471218 351598 471454
rect 351362 470898 351598 471134
rect 274562 453218 274798 453454
rect 274562 452898 274798 453134
rect 305282 453218 305518 453454
rect 305282 452898 305518 453134
rect 336002 453218 336238 453454
rect 336002 452898 336238 453134
rect 259202 435218 259438 435454
rect 259202 434898 259438 435134
rect 289922 435218 290158 435454
rect 289922 434898 290158 435134
rect 320642 435218 320878 435454
rect 320642 434898 320878 435134
rect 351362 435218 351598 435454
rect 351362 434898 351598 435134
rect 274562 417218 274798 417454
rect 274562 416898 274798 417134
rect 305282 417218 305518 417454
rect 305282 416898 305518 417134
rect 336002 417218 336238 417454
rect 336002 416898 336238 417134
rect 259202 399218 259438 399454
rect 259202 398898 259438 399134
rect 289922 399218 290158 399454
rect 289922 398898 290158 399134
rect 320642 399218 320878 399454
rect 320642 398898 320878 399134
rect 351362 399218 351598 399454
rect 351362 398898 351598 399134
rect 274562 381218 274798 381454
rect 274562 380898 274798 381134
rect 305282 381218 305518 381454
rect 305282 380898 305518 381134
rect 336002 381218 336238 381454
rect 336002 380898 336238 381134
rect 259202 363218 259438 363454
rect 259202 362898 259438 363134
rect 289922 363218 290158 363454
rect 289922 362898 290158 363134
rect 320642 363218 320878 363454
rect 320642 362898 320878 363134
rect 351362 363218 351598 363454
rect 351362 362898 351598 363134
rect 274562 345218 274798 345454
rect 274562 344898 274798 345134
rect 305282 345218 305518 345454
rect 305282 344898 305518 345134
rect 336002 345218 336238 345454
rect 336002 344898 336238 345134
rect 259202 327218 259438 327454
rect 259202 326898 259438 327134
rect 289922 327218 290158 327454
rect 289922 326898 290158 327134
rect 320642 327218 320878 327454
rect 320642 326898 320878 327134
rect 351362 327218 351598 327454
rect 351362 326898 351598 327134
rect 274562 309218 274798 309454
rect 274562 308898 274798 309134
rect 305282 309218 305518 309454
rect 305282 308898 305518 309134
rect 336002 309218 336238 309454
rect 336002 308898 336238 309134
rect 259202 291218 259438 291454
rect 259202 290898 259438 291134
rect 289922 291218 290158 291454
rect 289922 290898 290158 291134
rect 320642 291218 320878 291454
rect 320642 290898 320878 291134
rect 351362 291218 351598 291454
rect 351362 290898 351598 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 382082 687218 382318 687454
rect 382082 686898 382318 687134
rect 412802 687218 413038 687454
rect 412802 686898 413038 687134
rect 443522 687218 443758 687454
rect 443522 686898 443758 687134
rect 474242 687218 474478 687454
rect 474242 686898 474478 687134
rect 504962 687218 505198 687454
rect 504962 686898 505198 687134
rect 366722 669218 366958 669454
rect 366722 668898 366958 669134
rect 397442 669218 397678 669454
rect 397442 668898 397678 669134
rect 428162 669218 428398 669454
rect 428162 668898 428398 669134
rect 458882 669218 459118 669454
rect 458882 668898 459118 669134
rect 489602 669218 489838 669454
rect 489602 668898 489838 669134
rect 382082 651218 382318 651454
rect 382082 650898 382318 651134
rect 412802 651218 413038 651454
rect 412802 650898 413038 651134
rect 443522 651218 443758 651454
rect 443522 650898 443758 651134
rect 474242 651218 474478 651454
rect 474242 650898 474478 651134
rect 504962 651218 505198 651454
rect 504962 650898 505198 651134
rect 366722 633218 366958 633454
rect 366722 632898 366958 633134
rect 397442 633218 397678 633454
rect 397442 632898 397678 633134
rect 428162 633218 428398 633454
rect 428162 632898 428398 633134
rect 458882 633218 459118 633454
rect 458882 632898 459118 633134
rect 489602 633218 489838 633454
rect 489602 632898 489838 633134
rect 382082 615218 382318 615454
rect 382082 614898 382318 615134
rect 412802 615218 413038 615454
rect 412802 614898 413038 615134
rect 443522 615218 443758 615454
rect 443522 614898 443758 615134
rect 474242 615218 474478 615454
rect 474242 614898 474478 615134
rect 504962 615218 505198 615454
rect 504962 614898 505198 615134
rect 366722 597218 366958 597454
rect 366722 596898 366958 597134
rect 397442 597218 397678 597454
rect 397442 596898 397678 597134
rect 428162 597218 428398 597454
rect 428162 596898 428398 597134
rect 458882 597218 459118 597454
rect 458882 596898 459118 597134
rect 489602 597218 489838 597454
rect 489602 596898 489838 597134
rect 382082 579218 382318 579454
rect 382082 578898 382318 579134
rect 412802 579218 413038 579454
rect 412802 578898 413038 579134
rect 443522 579218 443758 579454
rect 443522 578898 443758 579134
rect 474242 579218 474478 579454
rect 474242 578898 474478 579134
rect 504962 579218 505198 579454
rect 504962 578898 505198 579134
rect 366722 561218 366958 561454
rect 366722 560898 366958 561134
rect 397442 561218 397678 561454
rect 397442 560898 397678 561134
rect 428162 561218 428398 561454
rect 428162 560898 428398 561134
rect 458882 561218 459118 561454
rect 458882 560898 459118 561134
rect 489602 561218 489838 561454
rect 489602 560898 489838 561134
rect 382082 543218 382318 543454
rect 382082 542898 382318 543134
rect 412802 543218 413038 543454
rect 412802 542898 413038 543134
rect 443522 543218 443758 543454
rect 443522 542898 443758 543134
rect 474242 543218 474478 543454
rect 474242 542898 474478 543134
rect 504962 543218 505198 543454
rect 504962 542898 505198 543134
rect 366722 525218 366958 525454
rect 366722 524898 366958 525134
rect 397442 525218 397678 525454
rect 397442 524898 397678 525134
rect 428162 525218 428398 525454
rect 428162 524898 428398 525134
rect 458882 525218 459118 525454
rect 458882 524898 459118 525134
rect 489602 525218 489838 525454
rect 489602 524898 489838 525134
rect 382082 507218 382318 507454
rect 382082 506898 382318 507134
rect 412802 507218 413038 507454
rect 412802 506898 413038 507134
rect 443522 507218 443758 507454
rect 443522 506898 443758 507134
rect 474242 507218 474478 507454
rect 474242 506898 474478 507134
rect 504962 507218 505198 507454
rect 504962 506898 505198 507134
rect 366722 489218 366958 489454
rect 366722 488898 366958 489134
rect 397442 489218 397678 489454
rect 397442 488898 397678 489134
rect 428162 489218 428398 489454
rect 428162 488898 428398 489134
rect 458882 489218 459118 489454
rect 458882 488898 459118 489134
rect 489602 489218 489838 489454
rect 489602 488898 489838 489134
rect 382082 471218 382318 471454
rect 382082 470898 382318 471134
rect 412802 471218 413038 471454
rect 412802 470898 413038 471134
rect 443522 471218 443758 471454
rect 443522 470898 443758 471134
rect 474242 471218 474478 471454
rect 474242 470898 474478 471134
rect 504962 471218 505198 471454
rect 504962 470898 505198 471134
rect 366722 453218 366958 453454
rect 366722 452898 366958 453134
rect 397442 453218 397678 453454
rect 397442 452898 397678 453134
rect 428162 453218 428398 453454
rect 428162 452898 428398 453134
rect 458882 453218 459118 453454
rect 458882 452898 459118 453134
rect 489602 453218 489838 453454
rect 489602 452898 489838 453134
rect 382082 435218 382318 435454
rect 382082 434898 382318 435134
rect 412802 435218 413038 435454
rect 412802 434898 413038 435134
rect 443522 435218 443758 435454
rect 443522 434898 443758 435134
rect 474242 435218 474478 435454
rect 474242 434898 474478 435134
rect 504962 435218 505198 435454
rect 504962 434898 505198 435134
rect 366722 417218 366958 417454
rect 366722 416898 366958 417134
rect 397442 417218 397678 417454
rect 397442 416898 397678 417134
rect 428162 417218 428398 417454
rect 428162 416898 428398 417134
rect 458882 417218 459118 417454
rect 458882 416898 459118 417134
rect 489602 417218 489838 417454
rect 489602 416898 489838 417134
rect 382082 399218 382318 399454
rect 382082 398898 382318 399134
rect 412802 399218 413038 399454
rect 412802 398898 413038 399134
rect 443522 399218 443758 399454
rect 443522 398898 443758 399134
rect 474242 399218 474478 399454
rect 474242 398898 474478 399134
rect 504962 399218 505198 399454
rect 504962 398898 505198 399134
rect 366722 381218 366958 381454
rect 366722 380898 366958 381134
rect 397442 381218 397678 381454
rect 397442 380898 397678 381134
rect 428162 381218 428398 381454
rect 428162 380898 428398 381134
rect 458882 381218 459118 381454
rect 458882 380898 459118 381134
rect 489602 381218 489838 381454
rect 489602 380898 489838 381134
rect 382082 363218 382318 363454
rect 382082 362898 382318 363134
rect 412802 363218 413038 363454
rect 412802 362898 413038 363134
rect 443522 363218 443758 363454
rect 443522 362898 443758 363134
rect 474242 363218 474478 363454
rect 474242 362898 474478 363134
rect 504962 363218 505198 363454
rect 504962 362898 505198 363134
rect 366722 345218 366958 345454
rect 366722 344898 366958 345134
rect 397442 345218 397678 345454
rect 397442 344898 397678 345134
rect 428162 345218 428398 345454
rect 428162 344898 428398 345134
rect 458882 345218 459118 345454
rect 458882 344898 459118 345134
rect 489602 345218 489838 345454
rect 489602 344898 489838 345134
rect 382082 327218 382318 327454
rect 382082 326898 382318 327134
rect 412802 327218 413038 327454
rect 412802 326898 413038 327134
rect 443522 327218 443758 327454
rect 443522 326898 443758 327134
rect 474242 327218 474478 327454
rect 474242 326898 474478 327134
rect 504962 327218 505198 327454
rect 504962 326898 505198 327134
rect 366722 309218 366958 309454
rect 366722 308898 366958 309134
rect 397442 309218 397678 309454
rect 397442 308898 397678 309134
rect 428162 309218 428398 309454
rect 428162 308898 428398 309134
rect 458882 309218 459118 309454
rect 458882 308898 459118 309134
rect 489602 309218 489838 309454
rect 489602 308898 489838 309134
rect 382082 291218 382318 291454
rect 382082 290898 382318 291134
rect 412802 291218 413038 291454
rect 412802 290898 413038 291134
rect 443522 291218 443758 291454
rect 443522 290898 443758 291134
rect 474242 291218 474478 291454
rect 474242 290898 474478 291134
rect 504962 291218 505198 291454
rect 504962 290898 505198 291134
rect 520322 669218 520558 669454
rect 520322 668898 520558 669134
rect 520322 633218 520558 633454
rect 520322 632898 520558 633134
rect 520322 597218 520558 597454
rect 520322 596898 520558 597134
rect 520322 561218 520558 561454
rect 520322 560898 520558 561134
rect 520322 525218 520558 525454
rect 520322 524898 520558 525134
rect 520322 489218 520558 489454
rect 520322 488898 520558 489134
rect 520322 453218 520558 453454
rect 520322 452898 520558 453134
rect 520322 417218 520558 417454
rect 520322 416898 520558 417134
rect 520322 381218 520558 381454
rect 520322 380898 520558 381134
rect 520322 345218 520558 345454
rect 520322 344898 520558 345134
rect 520322 309218 520558 309454
rect 520322 308898 520558 309134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 535682 687218 535918 687454
rect 535682 686898 535918 687134
rect 566402 687218 566638 687454
rect 566402 686898 566638 687134
rect 551042 669218 551278 669454
rect 551042 668898 551278 669134
rect 535682 651218 535918 651454
rect 535682 650898 535918 651134
rect 566402 651218 566638 651454
rect 566402 650898 566638 651134
rect 551042 633218 551278 633454
rect 551042 632898 551278 633134
rect 535682 615218 535918 615454
rect 535682 614898 535918 615134
rect 566402 615218 566638 615454
rect 566402 614898 566638 615134
rect 551042 597218 551278 597454
rect 551042 596898 551278 597134
rect 535682 579218 535918 579454
rect 535682 578898 535918 579134
rect 566402 579218 566638 579454
rect 566402 578898 566638 579134
rect 551042 561218 551278 561454
rect 551042 560898 551278 561134
rect 535682 543218 535918 543454
rect 535682 542898 535918 543134
rect 566402 543218 566638 543454
rect 566402 542898 566638 543134
rect 551042 525218 551278 525454
rect 551042 524898 551278 525134
rect 535682 507218 535918 507454
rect 535682 506898 535918 507134
rect 566402 507218 566638 507454
rect 566402 506898 566638 507134
rect 551042 489218 551278 489454
rect 551042 488898 551278 489134
rect 535682 471218 535918 471454
rect 535682 470898 535918 471134
rect 566402 471218 566638 471454
rect 566402 470898 566638 471134
rect 551042 453218 551278 453454
rect 551042 452898 551278 453134
rect 535682 435218 535918 435454
rect 535682 434898 535918 435134
rect 566402 435218 566638 435454
rect 566402 434898 566638 435134
rect 551042 417218 551278 417454
rect 551042 416898 551278 417134
rect 535682 399218 535918 399454
rect 535682 398898 535918 399134
rect 566402 399218 566638 399454
rect 566402 398898 566638 399134
rect 551042 381218 551278 381454
rect 551042 380898 551278 381134
rect 535682 363218 535918 363454
rect 535682 362898 535918 363134
rect 566402 363218 566638 363454
rect 566402 362898 566638 363134
rect 551042 345218 551278 345454
rect 551042 344898 551278 345134
rect 535682 327218 535918 327454
rect 535682 326898 535918 327134
rect 566402 327218 566638 327454
rect 566402 326898 566638 327134
rect 551042 309218 551278 309454
rect 551042 308898 551278 309134
rect 535682 291218 535918 291454
rect 535682 290898 535918 291134
rect 566402 291218 566638 291454
rect 566402 290898 566638 291134
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 167042 687454
rect 167278 687218 197762 687454
rect 197998 687218 228482 687454
rect 228718 687218 259202 687454
rect 259438 687218 289922 687454
rect 290158 687218 320642 687454
rect 320878 687218 351362 687454
rect 351598 687218 382082 687454
rect 382318 687218 412802 687454
rect 413038 687218 443522 687454
rect 443758 687218 474242 687454
rect 474478 687218 504962 687454
rect 505198 687218 535682 687454
rect 535918 687218 566402 687454
rect 566638 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 167042 687134
rect 167278 686898 197762 687134
rect 197998 686898 228482 687134
rect 228718 686898 259202 687134
rect 259438 686898 289922 687134
rect 290158 686898 320642 687134
rect 320878 686898 351362 687134
rect 351598 686898 382082 687134
rect 382318 686898 412802 687134
rect 413038 686898 443522 687134
rect 443758 686898 474242 687134
rect 474478 686898 504962 687134
rect 505198 686898 535682 687134
rect 535918 686898 566402 687134
rect 566638 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 182402 669454
rect 182638 669218 213122 669454
rect 213358 669218 243842 669454
rect 244078 669218 274562 669454
rect 274798 669218 305282 669454
rect 305518 669218 336002 669454
rect 336238 669218 366722 669454
rect 366958 669218 397442 669454
rect 397678 669218 428162 669454
rect 428398 669218 458882 669454
rect 459118 669218 489602 669454
rect 489838 669218 520322 669454
rect 520558 669218 551042 669454
rect 551278 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 182402 669134
rect 182638 668898 213122 669134
rect 213358 668898 243842 669134
rect 244078 668898 274562 669134
rect 274798 668898 305282 669134
rect 305518 668898 336002 669134
rect 336238 668898 366722 669134
rect 366958 668898 397442 669134
rect 397678 668898 428162 669134
rect 428398 668898 458882 669134
rect 459118 668898 489602 669134
rect 489838 668898 520322 669134
rect 520558 668898 551042 669134
rect 551278 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 167042 651454
rect 167278 651218 197762 651454
rect 197998 651218 228482 651454
rect 228718 651218 259202 651454
rect 259438 651218 289922 651454
rect 290158 651218 320642 651454
rect 320878 651218 351362 651454
rect 351598 651218 382082 651454
rect 382318 651218 412802 651454
rect 413038 651218 443522 651454
rect 443758 651218 474242 651454
rect 474478 651218 504962 651454
rect 505198 651218 535682 651454
rect 535918 651218 566402 651454
rect 566638 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 167042 651134
rect 167278 650898 197762 651134
rect 197998 650898 228482 651134
rect 228718 650898 259202 651134
rect 259438 650898 289922 651134
rect 290158 650898 320642 651134
rect 320878 650898 351362 651134
rect 351598 650898 382082 651134
rect 382318 650898 412802 651134
rect 413038 650898 443522 651134
rect 443758 650898 474242 651134
rect 474478 650898 504962 651134
rect 505198 650898 535682 651134
rect 535918 650898 566402 651134
rect 566638 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 182402 633454
rect 182638 633218 213122 633454
rect 213358 633218 243842 633454
rect 244078 633218 274562 633454
rect 274798 633218 305282 633454
rect 305518 633218 336002 633454
rect 336238 633218 366722 633454
rect 366958 633218 397442 633454
rect 397678 633218 428162 633454
rect 428398 633218 458882 633454
rect 459118 633218 489602 633454
rect 489838 633218 520322 633454
rect 520558 633218 551042 633454
rect 551278 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 182402 633134
rect 182638 632898 213122 633134
rect 213358 632898 243842 633134
rect 244078 632898 274562 633134
rect 274798 632898 305282 633134
rect 305518 632898 336002 633134
rect 336238 632898 366722 633134
rect 366958 632898 397442 633134
rect 397678 632898 428162 633134
rect 428398 632898 458882 633134
rect 459118 632898 489602 633134
rect 489838 632898 520322 633134
rect 520558 632898 551042 633134
rect 551278 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 167042 615454
rect 167278 615218 197762 615454
rect 197998 615218 228482 615454
rect 228718 615218 259202 615454
rect 259438 615218 289922 615454
rect 290158 615218 320642 615454
rect 320878 615218 351362 615454
rect 351598 615218 382082 615454
rect 382318 615218 412802 615454
rect 413038 615218 443522 615454
rect 443758 615218 474242 615454
rect 474478 615218 504962 615454
rect 505198 615218 535682 615454
rect 535918 615218 566402 615454
rect 566638 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 167042 615134
rect 167278 614898 197762 615134
rect 197998 614898 228482 615134
rect 228718 614898 259202 615134
rect 259438 614898 289922 615134
rect 290158 614898 320642 615134
rect 320878 614898 351362 615134
rect 351598 614898 382082 615134
rect 382318 614898 412802 615134
rect 413038 614898 443522 615134
rect 443758 614898 474242 615134
rect 474478 614898 504962 615134
rect 505198 614898 535682 615134
rect 535918 614898 566402 615134
rect 566638 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 182402 597454
rect 182638 597218 213122 597454
rect 213358 597218 243842 597454
rect 244078 597218 274562 597454
rect 274798 597218 305282 597454
rect 305518 597218 336002 597454
rect 336238 597218 366722 597454
rect 366958 597218 397442 597454
rect 397678 597218 428162 597454
rect 428398 597218 458882 597454
rect 459118 597218 489602 597454
rect 489838 597218 520322 597454
rect 520558 597218 551042 597454
rect 551278 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 182402 597134
rect 182638 596898 213122 597134
rect 213358 596898 243842 597134
rect 244078 596898 274562 597134
rect 274798 596898 305282 597134
rect 305518 596898 336002 597134
rect 336238 596898 366722 597134
rect 366958 596898 397442 597134
rect 397678 596898 428162 597134
rect 428398 596898 458882 597134
rect 459118 596898 489602 597134
rect 489838 596898 520322 597134
rect 520558 596898 551042 597134
rect 551278 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 167042 579454
rect 167278 579218 197762 579454
rect 197998 579218 228482 579454
rect 228718 579218 259202 579454
rect 259438 579218 289922 579454
rect 290158 579218 320642 579454
rect 320878 579218 351362 579454
rect 351598 579218 382082 579454
rect 382318 579218 412802 579454
rect 413038 579218 443522 579454
rect 443758 579218 474242 579454
rect 474478 579218 504962 579454
rect 505198 579218 535682 579454
rect 535918 579218 566402 579454
rect 566638 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 167042 579134
rect 167278 578898 197762 579134
rect 197998 578898 228482 579134
rect 228718 578898 259202 579134
rect 259438 578898 289922 579134
rect 290158 578898 320642 579134
rect 320878 578898 351362 579134
rect 351598 578898 382082 579134
rect 382318 578898 412802 579134
rect 413038 578898 443522 579134
rect 443758 578898 474242 579134
rect 474478 578898 504962 579134
rect 505198 578898 535682 579134
rect 535918 578898 566402 579134
rect 566638 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 182402 561454
rect 182638 561218 213122 561454
rect 213358 561218 243842 561454
rect 244078 561218 274562 561454
rect 274798 561218 305282 561454
rect 305518 561218 336002 561454
rect 336238 561218 366722 561454
rect 366958 561218 397442 561454
rect 397678 561218 428162 561454
rect 428398 561218 458882 561454
rect 459118 561218 489602 561454
rect 489838 561218 520322 561454
rect 520558 561218 551042 561454
rect 551278 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 182402 561134
rect 182638 560898 213122 561134
rect 213358 560898 243842 561134
rect 244078 560898 274562 561134
rect 274798 560898 305282 561134
rect 305518 560898 336002 561134
rect 336238 560898 366722 561134
rect 366958 560898 397442 561134
rect 397678 560898 428162 561134
rect 428398 560898 458882 561134
rect 459118 560898 489602 561134
rect 489838 560898 520322 561134
rect 520558 560898 551042 561134
rect 551278 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 167042 543454
rect 167278 543218 197762 543454
rect 197998 543218 228482 543454
rect 228718 543218 259202 543454
rect 259438 543218 289922 543454
rect 290158 543218 320642 543454
rect 320878 543218 351362 543454
rect 351598 543218 382082 543454
rect 382318 543218 412802 543454
rect 413038 543218 443522 543454
rect 443758 543218 474242 543454
rect 474478 543218 504962 543454
rect 505198 543218 535682 543454
rect 535918 543218 566402 543454
rect 566638 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 167042 543134
rect 167278 542898 197762 543134
rect 197998 542898 228482 543134
rect 228718 542898 259202 543134
rect 259438 542898 289922 543134
rect 290158 542898 320642 543134
rect 320878 542898 351362 543134
rect 351598 542898 382082 543134
rect 382318 542898 412802 543134
rect 413038 542898 443522 543134
rect 443758 542898 474242 543134
rect 474478 542898 504962 543134
rect 505198 542898 535682 543134
rect 535918 542898 566402 543134
rect 566638 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 182402 525454
rect 182638 525218 213122 525454
rect 213358 525218 243842 525454
rect 244078 525218 274562 525454
rect 274798 525218 305282 525454
rect 305518 525218 336002 525454
rect 336238 525218 366722 525454
rect 366958 525218 397442 525454
rect 397678 525218 428162 525454
rect 428398 525218 458882 525454
rect 459118 525218 489602 525454
rect 489838 525218 520322 525454
rect 520558 525218 551042 525454
rect 551278 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 182402 525134
rect 182638 524898 213122 525134
rect 213358 524898 243842 525134
rect 244078 524898 274562 525134
rect 274798 524898 305282 525134
rect 305518 524898 336002 525134
rect 336238 524898 366722 525134
rect 366958 524898 397442 525134
rect 397678 524898 428162 525134
rect 428398 524898 458882 525134
rect 459118 524898 489602 525134
rect 489838 524898 520322 525134
rect 520558 524898 551042 525134
rect 551278 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 167042 507454
rect 167278 507218 197762 507454
rect 197998 507218 228482 507454
rect 228718 507218 259202 507454
rect 259438 507218 289922 507454
rect 290158 507218 320642 507454
rect 320878 507218 351362 507454
rect 351598 507218 382082 507454
rect 382318 507218 412802 507454
rect 413038 507218 443522 507454
rect 443758 507218 474242 507454
rect 474478 507218 504962 507454
rect 505198 507218 535682 507454
rect 535918 507218 566402 507454
rect 566638 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 167042 507134
rect 167278 506898 197762 507134
rect 197998 506898 228482 507134
rect 228718 506898 259202 507134
rect 259438 506898 289922 507134
rect 290158 506898 320642 507134
rect 320878 506898 351362 507134
rect 351598 506898 382082 507134
rect 382318 506898 412802 507134
rect 413038 506898 443522 507134
rect 443758 506898 474242 507134
rect 474478 506898 504962 507134
rect 505198 506898 535682 507134
rect 535918 506898 566402 507134
rect 566638 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 182402 489454
rect 182638 489218 213122 489454
rect 213358 489218 243842 489454
rect 244078 489218 274562 489454
rect 274798 489218 305282 489454
rect 305518 489218 336002 489454
rect 336238 489218 366722 489454
rect 366958 489218 397442 489454
rect 397678 489218 428162 489454
rect 428398 489218 458882 489454
rect 459118 489218 489602 489454
rect 489838 489218 520322 489454
rect 520558 489218 551042 489454
rect 551278 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 182402 489134
rect 182638 488898 213122 489134
rect 213358 488898 243842 489134
rect 244078 488898 274562 489134
rect 274798 488898 305282 489134
rect 305518 488898 336002 489134
rect 336238 488898 366722 489134
rect 366958 488898 397442 489134
rect 397678 488898 428162 489134
rect 428398 488898 458882 489134
rect 459118 488898 489602 489134
rect 489838 488898 520322 489134
rect 520558 488898 551042 489134
rect 551278 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 167042 471454
rect 167278 471218 197762 471454
rect 197998 471218 228482 471454
rect 228718 471218 259202 471454
rect 259438 471218 289922 471454
rect 290158 471218 320642 471454
rect 320878 471218 351362 471454
rect 351598 471218 382082 471454
rect 382318 471218 412802 471454
rect 413038 471218 443522 471454
rect 443758 471218 474242 471454
rect 474478 471218 504962 471454
rect 505198 471218 535682 471454
rect 535918 471218 566402 471454
rect 566638 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 167042 471134
rect 167278 470898 197762 471134
rect 197998 470898 228482 471134
rect 228718 470898 259202 471134
rect 259438 470898 289922 471134
rect 290158 470898 320642 471134
rect 320878 470898 351362 471134
rect 351598 470898 382082 471134
rect 382318 470898 412802 471134
rect 413038 470898 443522 471134
rect 443758 470898 474242 471134
rect 474478 470898 504962 471134
rect 505198 470898 535682 471134
rect 535918 470898 566402 471134
rect 566638 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 182402 453454
rect 182638 453218 213122 453454
rect 213358 453218 243842 453454
rect 244078 453218 274562 453454
rect 274798 453218 305282 453454
rect 305518 453218 336002 453454
rect 336238 453218 366722 453454
rect 366958 453218 397442 453454
rect 397678 453218 428162 453454
rect 428398 453218 458882 453454
rect 459118 453218 489602 453454
rect 489838 453218 520322 453454
rect 520558 453218 551042 453454
rect 551278 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 182402 453134
rect 182638 452898 213122 453134
rect 213358 452898 243842 453134
rect 244078 452898 274562 453134
rect 274798 452898 305282 453134
rect 305518 452898 336002 453134
rect 336238 452898 366722 453134
rect 366958 452898 397442 453134
rect 397678 452898 428162 453134
rect 428398 452898 458882 453134
rect 459118 452898 489602 453134
rect 489838 452898 520322 453134
rect 520558 452898 551042 453134
rect 551278 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 167042 435454
rect 167278 435218 197762 435454
rect 197998 435218 228482 435454
rect 228718 435218 259202 435454
rect 259438 435218 289922 435454
rect 290158 435218 320642 435454
rect 320878 435218 351362 435454
rect 351598 435218 382082 435454
rect 382318 435218 412802 435454
rect 413038 435218 443522 435454
rect 443758 435218 474242 435454
rect 474478 435218 504962 435454
rect 505198 435218 535682 435454
rect 535918 435218 566402 435454
rect 566638 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 167042 435134
rect 167278 434898 197762 435134
rect 197998 434898 228482 435134
rect 228718 434898 259202 435134
rect 259438 434898 289922 435134
rect 290158 434898 320642 435134
rect 320878 434898 351362 435134
rect 351598 434898 382082 435134
rect 382318 434898 412802 435134
rect 413038 434898 443522 435134
rect 443758 434898 474242 435134
rect 474478 434898 504962 435134
rect 505198 434898 535682 435134
rect 535918 434898 566402 435134
rect 566638 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 182402 417454
rect 182638 417218 213122 417454
rect 213358 417218 243842 417454
rect 244078 417218 274562 417454
rect 274798 417218 305282 417454
rect 305518 417218 336002 417454
rect 336238 417218 366722 417454
rect 366958 417218 397442 417454
rect 397678 417218 428162 417454
rect 428398 417218 458882 417454
rect 459118 417218 489602 417454
rect 489838 417218 520322 417454
rect 520558 417218 551042 417454
rect 551278 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 182402 417134
rect 182638 416898 213122 417134
rect 213358 416898 243842 417134
rect 244078 416898 274562 417134
rect 274798 416898 305282 417134
rect 305518 416898 336002 417134
rect 336238 416898 366722 417134
rect 366958 416898 397442 417134
rect 397678 416898 428162 417134
rect 428398 416898 458882 417134
rect 459118 416898 489602 417134
rect 489838 416898 520322 417134
rect 520558 416898 551042 417134
rect 551278 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 167042 399454
rect 167278 399218 197762 399454
rect 197998 399218 228482 399454
rect 228718 399218 259202 399454
rect 259438 399218 289922 399454
rect 290158 399218 320642 399454
rect 320878 399218 351362 399454
rect 351598 399218 382082 399454
rect 382318 399218 412802 399454
rect 413038 399218 443522 399454
rect 443758 399218 474242 399454
rect 474478 399218 504962 399454
rect 505198 399218 535682 399454
rect 535918 399218 566402 399454
rect 566638 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 167042 399134
rect 167278 398898 197762 399134
rect 197998 398898 228482 399134
rect 228718 398898 259202 399134
rect 259438 398898 289922 399134
rect 290158 398898 320642 399134
rect 320878 398898 351362 399134
rect 351598 398898 382082 399134
rect 382318 398898 412802 399134
rect 413038 398898 443522 399134
rect 443758 398898 474242 399134
rect 474478 398898 504962 399134
rect 505198 398898 535682 399134
rect 535918 398898 566402 399134
rect 566638 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 182402 381454
rect 182638 381218 213122 381454
rect 213358 381218 243842 381454
rect 244078 381218 274562 381454
rect 274798 381218 305282 381454
rect 305518 381218 336002 381454
rect 336238 381218 366722 381454
rect 366958 381218 397442 381454
rect 397678 381218 428162 381454
rect 428398 381218 458882 381454
rect 459118 381218 489602 381454
rect 489838 381218 520322 381454
rect 520558 381218 551042 381454
rect 551278 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 182402 381134
rect 182638 380898 213122 381134
rect 213358 380898 243842 381134
rect 244078 380898 274562 381134
rect 274798 380898 305282 381134
rect 305518 380898 336002 381134
rect 336238 380898 366722 381134
rect 366958 380898 397442 381134
rect 397678 380898 428162 381134
rect 428398 380898 458882 381134
rect 459118 380898 489602 381134
rect 489838 380898 520322 381134
rect 520558 380898 551042 381134
rect 551278 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 167042 363454
rect 167278 363218 197762 363454
rect 197998 363218 228482 363454
rect 228718 363218 259202 363454
rect 259438 363218 289922 363454
rect 290158 363218 320642 363454
rect 320878 363218 351362 363454
rect 351598 363218 382082 363454
rect 382318 363218 412802 363454
rect 413038 363218 443522 363454
rect 443758 363218 474242 363454
rect 474478 363218 504962 363454
rect 505198 363218 535682 363454
rect 535918 363218 566402 363454
rect 566638 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 167042 363134
rect 167278 362898 197762 363134
rect 197998 362898 228482 363134
rect 228718 362898 259202 363134
rect 259438 362898 289922 363134
rect 290158 362898 320642 363134
rect 320878 362898 351362 363134
rect 351598 362898 382082 363134
rect 382318 362898 412802 363134
rect 413038 362898 443522 363134
rect 443758 362898 474242 363134
rect 474478 362898 504962 363134
rect 505198 362898 535682 363134
rect 535918 362898 566402 363134
rect 566638 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 182402 345454
rect 182638 345218 213122 345454
rect 213358 345218 243842 345454
rect 244078 345218 274562 345454
rect 274798 345218 305282 345454
rect 305518 345218 336002 345454
rect 336238 345218 366722 345454
rect 366958 345218 397442 345454
rect 397678 345218 428162 345454
rect 428398 345218 458882 345454
rect 459118 345218 489602 345454
rect 489838 345218 520322 345454
rect 520558 345218 551042 345454
rect 551278 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 182402 345134
rect 182638 344898 213122 345134
rect 213358 344898 243842 345134
rect 244078 344898 274562 345134
rect 274798 344898 305282 345134
rect 305518 344898 336002 345134
rect 336238 344898 366722 345134
rect 366958 344898 397442 345134
rect 397678 344898 428162 345134
rect 428398 344898 458882 345134
rect 459118 344898 489602 345134
rect 489838 344898 520322 345134
rect 520558 344898 551042 345134
rect 551278 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 167042 327454
rect 167278 327218 197762 327454
rect 197998 327218 228482 327454
rect 228718 327218 259202 327454
rect 259438 327218 289922 327454
rect 290158 327218 320642 327454
rect 320878 327218 351362 327454
rect 351598 327218 382082 327454
rect 382318 327218 412802 327454
rect 413038 327218 443522 327454
rect 443758 327218 474242 327454
rect 474478 327218 504962 327454
rect 505198 327218 535682 327454
rect 535918 327218 566402 327454
rect 566638 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 167042 327134
rect 167278 326898 197762 327134
rect 197998 326898 228482 327134
rect 228718 326898 259202 327134
rect 259438 326898 289922 327134
rect 290158 326898 320642 327134
rect 320878 326898 351362 327134
rect 351598 326898 382082 327134
rect 382318 326898 412802 327134
rect 413038 326898 443522 327134
rect 443758 326898 474242 327134
rect 474478 326898 504962 327134
rect 505198 326898 535682 327134
rect 535918 326898 566402 327134
rect 566638 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 182402 309454
rect 182638 309218 213122 309454
rect 213358 309218 243842 309454
rect 244078 309218 274562 309454
rect 274798 309218 305282 309454
rect 305518 309218 336002 309454
rect 336238 309218 366722 309454
rect 366958 309218 397442 309454
rect 397678 309218 428162 309454
rect 428398 309218 458882 309454
rect 459118 309218 489602 309454
rect 489838 309218 520322 309454
rect 520558 309218 551042 309454
rect 551278 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 182402 309134
rect 182638 308898 213122 309134
rect 213358 308898 243842 309134
rect 244078 308898 274562 309134
rect 274798 308898 305282 309134
rect 305518 308898 336002 309134
rect 336238 308898 366722 309134
rect 366958 308898 397442 309134
rect 397678 308898 428162 309134
rect 428398 308898 458882 309134
rect 459118 308898 489602 309134
rect 489838 308898 520322 309134
rect 520558 308898 551042 309134
rect 551278 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 167042 291454
rect 167278 291218 197762 291454
rect 197998 291218 228482 291454
rect 228718 291218 259202 291454
rect 259438 291218 289922 291454
rect 290158 291218 320642 291454
rect 320878 291218 351362 291454
rect 351598 291218 382082 291454
rect 382318 291218 412802 291454
rect 413038 291218 443522 291454
rect 443758 291218 474242 291454
rect 474478 291218 504962 291454
rect 505198 291218 535682 291454
rect 535918 291218 566402 291454
rect 566638 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 167042 291134
rect 167278 290898 197762 291134
rect 197998 290898 228482 291134
rect 228718 290898 259202 291134
rect 259438 290898 289922 291134
rect 290158 290898 320642 291134
rect 320878 290898 351362 291134
rect 351598 290898 382082 291134
rect 382318 290898 412802 291134
rect 413038 290898 443522 291134
rect 443758 290898 474242 291134
rect 474478 290898 504962 291134
rect 505198 290898 535682 291134
rect 535918 290898 566402 291134
rect 566638 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use computer  computer
timestamp 1635000722
transform 1 0 162792 0 1 281792
box 382 0 419506 420000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 281792 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 701792 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 701792 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 701792 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 701792 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 701792 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 701792 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 701792 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 701792 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 701792 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 701792 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 701792 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 701792 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 279792 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 703792 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 703792 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 703792 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 703792 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 703792 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 703792 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 703792 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 703792 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 703792 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 703792 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 703792 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 703792 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 279792 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 703792 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 703792 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 703792 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 703792 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 703792 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 703792 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 703792 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 703792 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 703792 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 703792 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 703792 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 279792 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 703792 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 703792 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 703792 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 703792 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 703792 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 703792 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 703792 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 703792 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 703792 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 703792 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 703792 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 279792 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 703792 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 703792 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 703792 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 703792 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 703792 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 703792 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 703792 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 703792 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 703792 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 703792 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 703792 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 703792 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 279792 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 703792 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 703792 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 703792 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 703792 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 703792 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 703792 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 703792 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 703792 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 703792 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 703792 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 703792 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 703792 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 281792 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 701792 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 701792 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 701792 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 701792 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 701792 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 701792 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 701792 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 701792 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 701792 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 701792 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 701792 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 701792 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 279792 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 703792 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 703792 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 703792 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 703792 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 703792 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 703792 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 703792 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 703792 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 703792 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 703792 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 703792 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 703792 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
