magic
tech sky130A
magscale 1 2
timestamp 1634858302
<< obsli1 >>
rect 1104 2159 459511 457521
<< obsm1 >>
rect 474 2128 459526 457552
<< metal2 >>
rect 1950 459200 2006 460000
rect 5906 459200 5962 460000
rect 9954 459200 10010 460000
rect 14002 459200 14058 460000
rect 18050 459200 18106 460000
rect 22098 459200 22154 460000
rect 26146 459200 26202 460000
rect 30194 459200 30250 460000
rect 34150 459200 34206 460000
rect 38198 459200 38254 460000
rect 42246 459200 42302 460000
rect 46294 459200 46350 460000
rect 50342 459200 50398 460000
rect 54390 459200 54446 460000
rect 58438 459200 58494 460000
rect 62394 459200 62450 460000
rect 66442 459200 66498 460000
rect 70490 459200 70546 460000
rect 74538 459200 74594 460000
rect 78586 459200 78642 460000
rect 82634 459200 82690 460000
rect 86682 459200 86738 460000
rect 90638 459200 90694 460000
rect 94686 459200 94742 460000
rect 98734 459200 98790 460000
rect 102782 459200 102838 460000
rect 106830 459200 106886 460000
rect 110878 459200 110934 460000
rect 114926 459200 114982 460000
rect 118882 459200 118938 460000
rect 122930 459200 122986 460000
rect 126978 459200 127034 460000
rect 131026 459200 131082 460000
rect 135074 459200 135130 460000
rect 139122 459200 139178 460000
rect 143170 459200 143226 460000
rect 147126 459200 147182 460000
rect 151174 459200 151230 460000
rect 155222 459200 155278 460000
rect 159270 459200 159326 460000
rect 163318 459200 163374 460000
rect 167366 459200 167422 460000
rect 171414 459200 171470 460000
rect 175370 459200 175426 460000
rect 179418 459200 179474 460000
rect 183466 459200 183522 460000
rect 187514 459200 187570 460000
rect 191562 459200 191618 460000
rect 195610 459200 195666 460000
rect 199658 459200 199714 460000
rect 203614 459200 203670 460000
rect 207662 459200 207718 460000
rect 211710 459200 211766 460000
rect 215758 459200 215814 460000
rect 219806 459200 219862 460000
rect 223854 459200 223910 460000
rect 227902 459200 227958 460000
rect 231950 459200 232006 460000
rect 235906 459200 235962 460000
rect 239954 459200 240010 460000
rect 244002 459200 244058 460000
rect 248050 459200 248106 460000
rect 252098 459200 252154 460000
rect 256146 459200 256202 460000
rect 260194 459200 260250 460000
rect 264150 459200 264206 460000
rect 268198 459200 268254 460000
rect 272246 459200 272302 460000
rect 276294 459200 276350 460000
rect 280342 459200 280398 460000
rect 284390 459200 284446 460000
rect 288438 459200 288494 460000
rect 292394 459200 292450 460000
rect 296442 459200 296498 460000
rect 300490 459200 300546 460000
rect 304538 459200 304594 460000
rect 308586 459200 308642 460000
rect 312634 459200 312690 460000
rect 316682 459200 316738 460000
rect 320638 459200 320694 460000
rect 324686 459200 324742 460000
rect 328734 459200 328790 460000
rect 332782 459200 332838 460000
rect 336830 459200 336886 460000
rect 340878 459200 340934 460000
rect 344926 459200 344982 460000
rect 348882 459200 348938 460000
rect 352930 459200 352986 460000
rect 356978 459200 357034 460000
rect 361026 459200 361082 460000
rect 365074 459200 365130 460000
rect 369122 459200 369178 460000
rect 373170 459200 373226 460000
rect 377126 459200 377182 460000
rect 381174 459200 381230 460000
rect 385222 459200 385278 460000
rect 389270 459200 389326 460000
rect 393318 459200 393374 460000
rect 397366 459200 397422 460000
rect 401414 459200 401470 460000
rect 405370 459200 405426 460000
rect 409418 459200 409474 460000
rect 413466 459200 413522 460000
rect 417514 459200 417570 460000
rect 421562 459200 421618 460000
rect 425610 459200 425666 460000
rect 429658 459200 429714 460000
rect 433614 459200 433670 460000
rect 437662 459200 437718 460000
rect 441710 459200 441766 460000
rect 445758 459200 445814 460000
rect 449806 459200 449862 460000
rect 453854 459200 453910 460000
rect 457902 459200 457958 460000
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 5078 0 5134 800
rect 5998 0 6054 800
rect 6918 0 6974 800
rect 7930 0 7986 800
rect 8850 0 8906 800
rect 9770 0 9826 800
rect 10690 0 10746 800
rect 11610 0 11666 800
rect 12530 0 12586 800
rect 13450 0 13506 800
rect 14462 0 14518 800
rect 15382 0 15438 800
rect 16302 0 16358 800
rect 17222 0 17278 800
rect 18142 0 18198 800
rect 19062 0 19118 800
rect 19982 0 20038 800
rect 20994 0 21050 800
rect 21914 0 21970 800
rect 22834 0 22890 800
rect 23754 0 23810 800
rect 24674 0 24730 800
rect 25594 0 25650 800
rect 26514 0 26570 800
rect 27526 0 27582 800
rect 28446 0 28502 800
rect 29366 0 29422 800
rect 30286 0 30342 800
rect 31206 0 31262 800
rect 32126 0 32182 800
rect 33046 0 33102 800
rect 34058 0 34114 800
rect 34978 0 35034 800
rect 35898 0 35954 800
rect 36818 0 36874 800
rect 37738 0 37794 800
rect 38658 0 38714 800
rect 39578 0 39634 800
rect 40590 0 40646 800
rect 41510 0 41566 800
rect 42430 0 42486 800
rect 43350 0 43406 800
rect 44270 0 44326 800
rect 45190 0 45246 800
rect 46110 0 46166 800
rect 47122 0 47178 800
rect 48042 0 48098 800
rect 48962 0 49018 800
rect 49882 0 49938 800
rect 50802 0 50858 800
rect 51722 0 51778 800
rect 52642 0 52698 800
rect 53654 0 53710 800
rect 54574 0 54630 800
rect 55494 0 55550 800
rect 56414 0 56470 800
rect 57334 0 57390 800
rect 58254 0 58310 800
rect 59174 0 59230 800
rect 60186 0 60242 800
rect 61106 0 61162 800
rect 62026 0 62082 800
rect 62946 0 63002 800
rect 63866 0 63922 800
rect 64786 0 64842 800
rect 65706 0 65762 800
rect 66718 0 66774 800
rect 67638 0 67694 800
rect 68558 0 68614 800
rect 69478 0 69534 800
rect 70398 0 70454 800
rect 71318 0 71374 800
rect 72238 0 72294 800
rect 73250 0 73306 800
rect 74170 0 74226 800
rect 75090 0 75146 800
rect 76010 0 76066 800
rect 76930 0 76986 800
rect 77850 0 77906 800
rect 78770 0 78826 800
rect 79782 0 79838 800
rect 80702 0 80758 800
rect 81622 0 81678 800
rect 82542 0 82598 800
rect 83462 0 83518 800
rect 84382 0 84438 800
rect 85302 0 85358 800
rect 86314 0 86370 800
rect 87234 0 87290 800
rect 88154 0 88210 800
rect 89074 0 89130 800
rect 89994 0 90050 800
rect 90914 0 90970 800
rect 91834 0 91890 800
rect 92846 0 92902 800
rect 93766 0 93822 800
rect 94686 0 94742 800
rect 95606 0 95662 800
rect 96526 0 96582 800
rect 97446 0 97502 800
rect 98366 0 98422 800
rect 99378 0 99434 800
rect 100298 0 100354 800
rect 101218 0 101274 800
rect 102138 0 102194 800
rect 103058 0 103114 800
rect 103978 0 104034 800
rect 104898 0 104954 800
rect 105910 0 105966 800
rect 106830 0 106886 800
rect 107750 0 107806 800
rect 108670 0 108726 800
rect 109590 0 109646 800
rect 110510 0 110566 800
rect 111430 0 111486 800
rect 112442 0 112498 800
rect 113362 0 113418 800
rect 114282 0 114338 800
rect 115202 0 115258 800
rect 116122 0 116178 800
rect 117042 0 117098 800
rect 117962 0 118018 800
rect 118974 0 119030 800
rect 119894 0 119950 800
rect 120814 0 120870 800
rect 121734 0 121790 800
rect 122654 0 122710 800
rect 123574 0 123630 800
rect 124494 0 124550 800
rect 125506 0 125562 800
rect 126426 0 126482 800
rect 127346 0 127402 800
rect 128266 0 128322 800
rect 129186 0 129242 800
rect 130106 0 130162 800
rect 131026 0 131082 800
rect 132038 0 132094 800
rect 132958 0 133014 800
rect 133878 0 133934 800
rect 134798 0 134854 800
rect 135718 0 135774 800
rect 136638 0 136694 800
rect 137558 0 137614 800
rect 138570 0 138626 800
rect 139490 0 139546 800
rect 140410 0 140466 800
rect 141330 0 141386 800
rect 142250 0 142306 800
rect 143170 0 143226 800
rect 144090 0 144146 800
rect 145102 0 145158 800
rect 146022 0 146078 800
rect 146942 0 146998 800
rect 147862 0 147918 800
rect 148782 0 148838 800
rect 149702 0 149758 800
rect 150622 0 150678 800
rect 151634 0 151690 800
rect 152554 0 152610 800
rect 153474 0 153530 800
rect 154394 0 154450 800
rect 155314 0 155370 800
rect 156234 0 156290 800
rect 157154 0 157210 800
rect 158074 0 158130 800
rect 159086 0 159142 800
rect 160006 0 160062 800
rect 160926 0 160982 800
rect 161846 0 161902 800
rect 162766 0 162822 800
rect 163686 0 163742 800
rect 164606 0 164662 800
rect 165618 0 165674 800
rect 166538 0 166594 800
rect 167458 0 167514 800
rect 168378 0 168434 800
rect 169298 0 169354 800
rect 170218 0 170274 800
rect 171138 0 171194 800
rect 172150 0 172206 800
rect 173070 0 173126 800
rect 173990 0 174046 800
rect 174910 0 174966 800
rect 175830 0 175886 800
rect 176750 0 176806 800
rect 177670 0 177726 800
rect 178682 0 178738 800
rect 179602 0 179658 800
rect 180522 0 180578 800
rect 181442 0 181498 800
rect 182362 0 182418 800
rect 183282 0 183338 800
rect 184202 0 184258 800
rect 185214 0 185270 800
rect 186134 0 186190 800
rect 187054 0 187110 800
rect 187974 0 188030 800
rect 188894 0 188950 800
rect 189814 0 189870 800
rect 190734 0 190790 800
rect 191746 0 191802 800
rect 192666 0 192722 800
rect 193586 0 193642 800
rect 194506 0 194562 800
rect 195426 0 195482 800
rect 196346 0 196402 800
rect 197266 0 197322 800
rect 198278 0 198334 800
rect 199198 0 199254 800
rect 200118 0 200174 800
rect 201038 0 201094 800
rect 201958 0 202014 800
rect 202878 0 202934 800
rect 203798 0 203854 800
rect 204810 0 204866 800
rect 205730 0 205786 800
rect 206650 0 206706 800
rect 207570 0 207626 800
rect 208490 0 208546 800
rect 209410 0 209466 800
rect 210330 0 210386 800
rect 211342 0 211398 800
rect 212262 0 212318 800
rect 213182 0 213238 800
rect 214102 0 214158 800
rect 215022 0 215078 800
rect 215942 0 215998 800
rect 216862 0 216918 800
rect 217874 0 217930 800
rect 218794 0 218850 800
rect 219714 0 219770 800
rect 220634 0 220690 800
rect 221554 0 221610 800
rect 222474 0 222530 800
rect 223394 0 223450 800
rect 224406 0 224462 800
rect 225326 0 225382 800
rect 226246 0 226302 800
rect 227166 0 227222 800
rect 228086 0 228142 800
rect 229006 0 229062 800
rect 229926 0 229982 800
rect 230938 0 230994 800
rect 231858 0 231914 800
rect 232778 0 232834 800
rect 233698 0 233754 800
rect 234618 0 234674 800
rect 235538 0 235594 800
rect 236458 0 236514 800
rect 237470 0 237526 800
rect 238390 0 238446 800
rect 239310 0 239366 800
rect 240230 0 240286 800
rect 241150 0 241206 800
rect 242070 0 242126 800
rect 242990 0 243046 800
rect 244002 0 244058 800
rect 244922 0 244978 800
rect 245842 0 245898 800
rect 246762 0 246818 800
rect 247682 0 247738 800
rect 248602 0 248658 800
rect 249522 0 249578 800
rect 250534 0 250590 800
rect 251454 0 251510 800
rect 252374 0 252430 800
rect 253294 0 253350 800
rect 254214 0 254270 800
rect 255134 0 255190 800
rect 256054 0 256110 800
rect 257066 0 257122 800
rect 257986 0 258042 800
rect 258906 0 258962 800
rect 259826 0 259882 800
rect 260746 0 260802 800
rect 261666 0 261722 800
rect 262586 0 262642 800
rect 263598 0 263654 800
rect 264518 0 264574 800
rect 265438 0 265494 800
rect 266358 0 266414 800
rect 267278 0 267334 800
rect 268198 0 268254 800
rect 269118 0 269174 800
rect 270130 0 270186 800
rect 271050 0 271106 800
rect 271970 0 272026 800
rect 272890 0 272946 800
rect 273810 0 273866 800
rect 274730 0 274786 800
rect 275650 0 275706 800
rect 276662 0 276718 800
rect 277582 0 277638 800
rect 278502 0 278558 800
rect 279422 0 279478 800
rect 280342 0 280398 800
rect 281262 0 281318 800
rect 282182 0 282238 800
rect 283194 0 283250 800
rect 284114 0 284170 800
rect 285034 0 285090 800
rect 285954 0 286010 800
rect 286874 0 286930 800
rect 287794 0 287850 800
rect 288714 0 288770 800
rect 289726 0 289782 800
rect 290646 0 290702 800
rect 291566 0 291622 800
rect 292486 0 292542 800
rect 293406 0 293462 800
rect 294326 0 294382 800
rect 295246 0 295302 800
rect 296258 0 296314 800
rect 297178 0 297234 800
rect 298098 0 298154 800
rect 299018 0 299074 800
rect 299938 0 299994 800
rect 300858 0 300914 800
rect 301778 0 301834 800
rect 302790 0 302846 800
rect 303710 0 303766 800
rect 304630 0 304686 800
rect 305550 0 305606 800
rect 306470 0 306526 800
rect 307390 0 307446 800
rect 308310 0 308366 800
rect 309230 0 309286 800
rect 310242 0 310298 800
rect 311162 0 311218 800
rect 312082 0 312138 800
rect 313002 0 313058 800
rect 313922 0 313978 800
rect 314842 0 314898 800
rect 315762 0 315818 800
rect 316774 0 316830 800
rect 317694 0 317750 800
rect 318614 0 318670 800
rect 319534 0 319590 800
rect 320454 0 320510 800
rect 321374 0 321430 800
rect 322294 0 322350 800
rect 323306 0 323362 800
rect 324226 0 324282 800
rect 325146 0 325202 800
rect 326066 0 326122 800
rect 326986 0 327042 800
rect 327906 0 327962 800
rect 328826 0 328882 800
rect 329838 0 329894 800
rect 330758 0 330814 800
rect 331678 0 331734 800
rect 332598 0 332654 800
rect 333518 0 333574 800
rect 334438 0 334494 800
rect 335358 0 335414 800
rect 336370 0 336426 800
rect 337290 0 337346 800
rect 338210 0 338266 800
rect 339130 0 339186 800
rect 340050 0 340106 800
rect 340970 0 341026 800
rect 341890 0 341946 800
rect 342902 0 342958 800
rect 343822 0 343878 800
rect 344742 0 344798 800
rect 345662 0 345718 800
rect 346582 0 346638 800
rect 347502 0 347558 800
rect 348422 0 348478 800
rect 349434 0 349490 800
rect 350354 0 350410 800
rect 351274 0 351330 800
rect 352194 0 352250 800
rect 353114 0 353170 800
rect 354034 0 354090 800
rect 354954 0 355010 800
rect 355966 0 356022 800
rect 356886 0 356942 800
rect 357806 0 357862 800
rect 358726 0 358782 800
rect 359646 0 359702 800
rect 360566 0 360622 800
rect 361486 0 361542 800
rect 362498 0 362554 800
rect 363418 0 363474 800
rect 364338 0 364394 800
rect 365258 0 365314 800
rect 366178 0 366234 800
rect 367098 0 367154 800
rect 368018 0 368074 800
rect 369030 0 369086 800
rect 369950 0 370006 800
rect 370870 0 370926 800
rect 371790 0 371846 800
rect 372710 0 372766 800
rect 373630 0 373686 800
rect 374550 0 374606 800
rect 375562 0 375618 800
rect 376482 0 376538 800
rect 377402 0 377458 800
rect 378322 0 378378 800
rect 379242 0 379298 800
rect 380162 0 380218 800
rect 381082 0 381138 800
rect 382094 0 382150 800
rect 383014 0 383070 800
rect 383934 0 383990 800
rect 384854 0 384910 800
rect 385774 0 385830 800
rect 386694 0 386750 800
rect 387614 0 387670 800
rect 388626 0 388682 800
rect 389546 0 389602 800
rect 390466 0 390522 800
rect 391386 0 391442 800
rect 392306 0 392362 800
rect 393226 0 393282 800
rect 394146 0 394202 800
rect 395158 0 395214 800
rect 396078 0 396134 800
rect 396998 0 397054 800
rect 397918 0 397974 800
rect 398838 0 398894 800
rect 399758 0 399814 800
rect 400678 0 400734 800
rect 401690 0 401746 800
rect 402610 0 402666 800
rect 403530 0 403586 800
rect 404450 0 404506 800
rect 405370 0 405426 800
rect 406290 0 406346 800
rect 407210 0 407266 800
rect 408222 0 408278 800
rect 409142 0 409198 800
rect 410062 0 410118 800
rect 410982 0 411038 800
rect 411902 0 411958 800
rect 412822 0 412878 800
rect 413742 0 413798 800
rect 414754 0 414810 800
rect 415674 0 415730 800
rect 416594 0 416650 800
rect 417514 0 417570 800
rect 418434 0 418490 800
rect 419354 0 419410 800
rect 420274 0 420330 800
rect 421286 0 421342 800
rect 422206 0 422262 800
rect 423126 0 423182 800
rect 424046 0 424102 800
rect 424966 0 425022 800
rect 425886 0 425942 800
rect 426806 0 426862 800
rect 427818 0 427874 800
rect 428738 0 428794 800
rect 429658 0 429714 800
rect 430578 0 430634 800
rect 431498 0 431554 800
rect 432418 0 432474 800
rect 433338 0 433394 800
rect 434350 0 434406 800
rect 435270 0 435326 800
rect 436190 0 436246 800
rect 437110 0 437166 800
rect 438030 0 438086 800
rect 438950 0 439006 800
rect 439870 0 439926 800
rect 440882 0 440938 800
rect 441802 0 441858 800
rect 442722 0 442778 800
rect 443642 0 443698 800
rect 444562 0 444618 800
rect 445482 0 445538 800
rect 446402 0 446458 800
rect 447414 0 447470 800
rect 448334 0 448390 800
rect 449254 0 449310 800
rect 450174 0 450230 800
rect 451094 0 451150 800
rect 452014 0 452070 800
rect 452934 0 452990 800
rect 453946 0 454002 800
rect 454866 0 454922 800
rect 455786 0 455842 800
rect 456706 0 456762 800
rect 457626 0 457682 800
rect 458546 0 458602 800
rect 459466 0 459522 800
<< obsm2 >>
rect 480 459144 1894 459218
rect 2062 459144 5850 459218
rect 6018 459144 9898 459218
rect 10066 459144 13946 459218
rect 14114 459144 17994 459218
rect 18162 459144 22042 459218
rect 22210 459144 26090 459218
rect 26258 459144 30138 459218
rect 30306 459144 34094 459218
rect 34262 459144 38142 459218
rect 38310 459144 42190 459218
rect 42358 459144 46238 459218
rect 46406 459144 50286 459218
rect 50454 459144 54334 459218
rect 54502 459144 58382 459218
rect 58550 459144 62338 459218
rect 62506 459144 66386 459218
rect 66554 459144 70434 459218
rect 70602 459144 74482 459218
rect 74650 459144 78530 459218
rect 78698 459144 82578 459218
rect 82746 459144 86626 459218
rect 86794 459144 90582 459218
rect 90750 459144 94630 459218
rect 94798 459144 98678 459218
rect 98846 459144 102726 459218
rect 102894 459144 106774 459218
rect 106942 459144 110822 459218
rect 110990 459144 114870 459218
rect 115038 459144 118826 459218
rect 118994 459144 122874 459218
rect 123042 459144 126922 459218
rect 127090 459144 130970 459218
rect 131138 459144 135018 459218
rect 135186 459144 139066 459218
rect 139234 459144 143114 459218
rect 143282 459144 147070 459218
rect 147238 459144 151118 459218
rect 151286 459144 155166 459218
rect 155334 459144 159214 459218
rect 159382 459144 163262 459218
rect 163430 459144 167310 459218
rect 167478 459144 171358 459218
rect 171526 459144 175314 459218
rect 175482 459144 179362 459218
rect 179530 459144 183410 459218
rect 183578 459144 187458 459218
rect 187626 459144 191506 459218
rect 191674 459144 195554 459218
rect 195722 459144 199602 459218
rect 199770 459144 203558 459218
rect 203726 459144 207606 459218
rect 207774 459144 211654 459218
rect 211822 459144 215702 459218
rect 215870 459144 219750 459218
rect 219918 459144 223798 459218
rect 223966 459144 227846 459218
rect 228014 459144 231894 459218
rect 232062 459144 235850 459218
rect 236018 459144 239898 459218
rect 240066 459144 243946 459218
rect 244114 459144 247994 459218
rect 248162 459144 252042 459218
rect 252210 459144 256090 459218
rect 256258 459144 260138 459218
rect 260306 459144 264094 459218
rect 264262 459144 268142 459218
rect 268310 459144 272190 459218
rect 272358 459144 276238 459218
rect 276406 459144 280286 459218
rect 280454 459144 284334 459218
rect 284502 459144 288382 459218
rect 288550 459144 292338 459218
rect 292506 459144 296386 459218
rect 296554 459144 300434 459218
rect 300602 459144 304482 459218
rect 304650 459144 308530 459218
rect 308698 459144 312578 459218
rect 312746 459144 316626 459218
rect 316794 459144 320582 459218
rect 320750 459144 324630 459218
rect 324798 459144 328678 459218
rect 328846 459144 332726 459218
rect 332894 459144 336774 459218
rect 336942 459144 340822 459218
rect 340990 459144 344870 459218
rect 345038 459144 348826 459218
rect 348994 459144 352874 459218
rect 353042 459144 356922 459218
rect 357090 459144 360970 459218
rect 361138 459144 365018 459218
rect 365186 459144 369066 459218
rect 369234 459144 373114 459218
rect 373282 459144 377070 459218
rect 377238 459144 381118 459218
rect 381286 459144 385166 459218
rect 385334 459144 389214 459218
rect 389382 459144 393262 459218
rect 393430 459144 397310 459218
rect 397478 459144 401358 459218
rect 401526 459144 405314 459218
rect 405482 459144 409362 459218
rect 409530 459144 413410 459218
rect 413578 459144 417458 459218
rect 417626 459144 421506 459218
rect 421674 459144 425554 459218
rect 425722 459144 429602 459218
rect 429770 459144 433558 459218
rect 433726 459144 437606 459218
rect 437774 459144 441654 459218
rect 441822 459144 445702 459218
rect 445870 459144 449750 459218
rect 449918 459144 453798 459218
rect 453966 459144 457846 459218
rect 458014 459144 459520 459218
rect 480 856 459520 459144
rect 590 734 1342 856
rect 1510 734 2262 856
rect 2430 734 3182 856
rect 3350 734 4102 856
rect 4270 734 5022 856
rect 5190 734 5942 856
rect 6110 734 6862 856
rect 7030 734 7874 856
rect 8042 734 8794 856
rect 8962 734 9714 856
rect 9882 734 10634 856
rect 10802 734 11554 856
rect 11722 734 12474 856
rect 12642 734 13394 856
rect 13562 734 14406 856
rect 14574 734 15326 856
rect 15494 734 16246 856
rect 16414 734 17166 856
rect 17334 734 18086 856
rect 18254 734 19006 856
rect 19174 734 19926 856
rect 20094 734 20938 856
rect 21106 734 21858 856
rect 22026 734 22778 856
rect 22946 734 23698 856
rect 23866 734 24618 856
rect 24786 734 25538 856
rect 25706 734 26458 856
rect 26626 734 27470 856
rect 27638 734 28390 856
rect 28558 734 29310 856
rect 29478 734 30230 856
rect 30398 734 31150 856
rect 31318 734 32070 856
rect 32238 734 32990 856
rect 33158 734 34002 856
rect 34170 734 34922 856
rect 35090 734 35842 856
rect 36010 734 36762 856
rect 36930 734 37682 856
rect 37850 734 38602 856
rect 38770 734 39522 856
rect 39690 734 40534 856
rect 40702 734 41454 856
rect 41622 734 42374 856
rect 42542 734 43294 856
rect 43462 734 44214 856
rect 44382 734 45134 856
rect 45302 734 46054 856
rect 46222 734 47066 856
rect 47234 734 47986 856
rect 48154 734 48906 856
rect 49074 734 49826 856
rect 49994 734 50746 856
rect 50914 734 51666 856
rect 51834 734 52586 856
rect 52754 734 53598 856
rect 53766 734 54518 856
rect 54686 734 55438 856
rect 55606 734 56358 856
rect 56526 734 57278 856
rect 57446 734 58198 856
rect 58366 734 59118 856
rect 59286 734 60130 856
rect 60298 734 61050 856
rect 61218 734 61970 856
rect 62138 734 62890 856
rect 63058 734 63810 856
rect 63978 734 64730 856
rect 64898 734 65650 856
rect 65818 734 66662 856
rect 66830 734 67582 856
rect 67750 734 68502 856
rect 68670 734 69422 856
rect 69590 734 70342 856
rect 70510 734 71262 856
rect 71430 734 72182 856
rect 72350 734 73194 856
rect 73362 734 74114 856
rect 74282 734 75034 856
rect 75202 734 75954 856
rect 76122 734 76874 856
rect 77042 734 77794 856
rect 77962 734 78714 856
rect 78882 734 79726 856
rect 79894 734 80646 856
rect 80814 734 81566 856
rect 81734 734 82486 856
rect 82654 734 83406 856
rect 83574 734 84326 856
rect 84494 734 85246 856
rect 85414 734 86258 856
rect 86426 734 87178 856
rect 87346 734 88098 856
rect 88266 734 89018 856
rect 89186 734 89938 856
rect 90106 734 90858 856
rect 91026 734 91778 856
rect 91946 734 92790 856
rect 92958 734 93710 856
rect 93878 734 94630 856
rect 94798 734 95550 856
rect 95718 734 96470 856
rect 96638 734 97390 856
rect 97558 734 98310 856
rect 98478 734 99322 856
rect 99490 734 100242 856
rect 100410 734 101162 856
rect 101330 734 102082 856
rect 102250 734 103002 856
rect 103170 734 103922 856
rect 104090 734 104842 856
rect 105010 734 105854 856
rect 106022 734 106774 856
rect 106942 734 107694 856
rect 107862 734 108614 856
rect 108782 734 109534 856
rect 109702 734 110454 856
rect 110622 734 111374 856
rect 111542 734 112386 856
rect 112554 734 113306 856
rect 113474 734 114226 856
rect 114394 734 115146 856
rect 115314 734 116066 856
rect 116234 734 116986 856
rect 117154 734 117906 856
rect 118074 734 118918 856
rect 119086 734 119838 856
rect 120006 734 120758 856
rect 120926 734 121678 856
rect 121846 734 122598 856
rect 122766 734 123518 856
rect 123686 734 124438 856
rect 124606 734 125450 856
rect 125618 734 126370 856
rect 126538 734 127290 856
rect 127458 734 128210 856
rect 128378 734 129130 856
rect 129298 734 130050 856
rect 130218 734 130970 856
rect 131138 734 131982 856
rect 132150 734 132902 856
rect 133070 734 133822 856
rect 133990 734 134742 856
rect 134910 734 135662 856
rect 135830 734 136582 856
rect 136750 734 137502 856
rect 137670 734 138514 856
rect 138682 734 139434 856
rect 139602 734 140354 856
rect 140522 734 141274 856
rect 141442 734 142194 856
rect 142362 734 143114 856
rect 143282 734 144034 856
rect 144202 734 145046 856
rect 145214 734 145966 856
rect 146134 734 146886 856
rect 147054 734 147806 856
rect 147974 734 148726 856
rect 148894 734 149646 856
rect 149814 734 150566 856
rect 150734 734 151578 856
rect 151746 734 152498 856
rect 152666 734 153418 856
rect 153586 734 154338 856
rect 154506 734 155258 856
rect 155426 734 156178 856
rect 156346 734 157098 856
rect 157266 734 158018 856
rect 158186 734 159030 856
rect 159198 734 159950 856
rect 160118 734 160870 856
rect 161038 734 161790 856
rect 161958 734 162710 856
rect 162878 734 163630 856
rect 163798 734 164550 856
rect 164718 734 165562 856
rect 165730 734 166482 856
rect 166650 734 167402 856
rect 167570 734 168322 856
rect 168490 734 169242 856
rect 169410 734 170162 856
rect 170330 734 171082 856
rect 171250 734 172094 856
rect 172262 734 173014 856
rect 173182 734 173934 856
rect 174102 734 174854 856
rect 175022 734 175774 856
rect 175942 734 176694 856
rect 176862 734 177614 856
rect 177782 734 178626 856
rect 178794 734 179546 856
rect 179714 734 180466 856
rect 180634 734 181386 856
rect 181554 734 182306 856
rect 182474 734 183226 856
rect 183394 734 184146 856
rect 184314 734 185158 856
rect 185326 734 186078 856
rect 186246 734 186998 856
rect 187166 734 187918 856
rect 188086 734 188838 856
rect 189006 734 189758 856
rect 189926 734 190678 856
rect 190846 734 191690 856
rect 191858 734 192610 856
rect 192778 734 193530 856
rect 193698 734 194450 856
rect 194618 734 195370 856
rect 195538 734 196290 856
rect 196458 734 197210 856
rect 197378 734 198222 856
rect 198390 734 199142 856
rect 199310 734 200062 856
rect 200230 734 200982 856
rect 201150 734 201902 856
rect 202070 734 202822 856
rect 202990 734 203742 856
rect 203910 734 204754 856
rect 204922 734 205674 856
rect 205842 734 206594 856
rect 206762 734 207514 856
rect 207682 734 208434 856
rect 208602 734 209354 856
rect 209522 734 210274 856
rect 210442 734 211286 856
rect 211454 734 212206 856
rect 212374 734 213126 856
rect 213294 734 214046 856
rect 214214 734 214966 856
rect 215134 734 215886 856
rect 216054 734 216806 856
rect 216974 734 217818 856
rect 217986 734 218738 856
rect 218906 734 219658 856
rect 219826 734 220578 856
rect 220746 734 221498 856
rect 221666 734 222418 856
rect 222586 734 223338 856
rect 223506 734 224350 856
rect 224518 734 225270 856
rect 225438 734 226190 856
rect 226358 734 227110 856
rect 227278 734 228030 856
rect 228198 734 228950 856
rect 229118 734 229870 856
rect 230038 734 230882 856
rect 231050 734 231802 856
rect 231970 734 232722 856
rect 232890 734 233642 856
rect 233810 734 234562 856
rect 234730 734 235482 856
rect 235650 734 236402 856
rect 236570 734 237414 856
rect 237582 734 238334 856
rect 238502 734 239254 856
rect 239422 734 240174 856
rect 240342 734 241094 856
rect 241262 734 242014 856
rect 242182 734 242934 856
rect 243102 734 243946 856
rect 244114 734 244866 856
rect 245034 734 245786 856
rect 245954 734 246706 856
rect 246874 734 247626 856
rect 247794 734 248546 856
rect 248714 734 249466 856
rect 249634 734 250478 856
rect 250646 734 251398 856
rect 251566 734 252318 856
rect 252486 734 253238 856
rect 253406 734 254158 856
rect 254326 734 255078 856
rect 255246 734 255998 856
rect 256166 734 257010 856
rect 257178 734 257930 856
rect 258098 734 258850 856
rect 259018 734 259770 856
rect 259938 734 260690 856
rect 260858 734 261610 856
rect 261778 734 262530 856
rect 262698 734 263542 856
rect 263710 734 264462 856
rect 264630 734 265382 856
rect 265550 734 266302 856
rect 266470 734 267222 856
rect 267390 734 268142 856
rect 268310 734 269062 856
rect 269230 734 270074 856
rect 270242 734 270994 856
rect 271162 734 271914 856
rect 272082 734 272834 856
rect 273002 734 273754 856
rect 273922 734 274674 856
rect 274842 734 275594 856
rect 275762 734 276606 856
rect 276774 734 277526 856
rect 277694 734 278446 856
rect 278614 734 279366 856
rect 279534 734 280286 856
rect 280454 734 281206 856
rect 281374 734 282126 856
rect 282294 734 283138 856
rect 283306 734 284058 856
rect 284226 734 284978 856
rect 285146 734 285898 856
rect 286066 734 286818 856
rect 286986 734 287738 856
rect 287906 734 288658 856
rect 288826 734 289670 856
rect 289838 734 290590 856
rect 290758 734 291510 856
rect 291678 734 292430 856
rect 292598 734 293350 856
rect 293518 734 294270 856
rect 294438 734 295190 856
rect 295358 734 296202 856
rect 296370 734 297122 856
rect 297290 734 298042 856
rect 298210 734 298962 856
rect 299130 734 299882 856
rect 300050 734 300802 856
rect 300970 734 301722 856
rect 301890 734 302734 856
rect 302902 734 303654 856
rect 303822 734 304574 856
rect 304742 734 305494 856
rect 305662 734 306414 856
rect 306582 734 307334 856
rect 307502 734 308254 856
rect 308422 734 309174 856
rect 309342 734 310186 856
rect 310354 734 311106 856
rect 311274 734 312026 856
rect 312194 734 312946 856
rect 313114 734 313866 856
rect 314034 734 314786 856
rect 314954 734 315706 856
rect 315874 734 316718 856
rect 316886 734 317638 856
rect 317806 734 318558 856
rect 318726 734 319478 856
rect 319646 734 320398 856
rect 320566 734 321318 856
rect 321486 734 322238 856
rect 322406 734 323250 856
rect 323418 734 324170 856
rect 324338 734 325090 856
rect 325258 734 326010 856
rect 326178 734 326930 856
rect 327098 734 327850 856
rect 328018 734 328770 856
rect 328938 734 329782 856
rect 329950 734 330702 856
rect 330870 734 331622 856
rect 331790 734 332542 856
rect 332710 734 333462 856
rect 333630 734 334382 856
rect 334550 734 335302 856
rect 335470 734 336314 856
rect 336482 734 337234 856
rect 337402 734 338154 856
rect 338322 734 339074 856
rect 339242 734 339994 856
rect 340162 734 340914 856
rect 341082 734 341834 856
rect 342002 734 342846 856
rect 343014 734 343766 856
rect 343934 734 344686 856
rect 344854 734 345606 856
rect 345774 734 346526 856
rect 346694 734 347446 856
rect 347614 734 348366 856
rect 348534 734 349378 856
rect 349546 734 350298 856
rect 350466 734 351218 856
rect 351386 734 352138 856
rect 352306 734 353058 856
rect 353226 734 353978 856
rect 354146 734 354898 856
rect 355066 734 355910 856
rect 356078 734 356830 856
rect 356998 734 357750 856
rect 357918 734 358670 856
rect 358838 734 359590 856
rect 359758 734 360510 856
rect 360678 734 361430 856
rect 361598 734 362442 856
rect 362610 734 363362 856
rect 363530 734 364282 856
rect 364450 734 365202 856
rect 365370 734 366122 856
rect 366290 734 367042 856
rect 367210 734 367962 856
rect 368130 734 368974 856
rect 369142 734 369894 856
rect 370062 734 370814 856
rect 370982 734 371734 856
rect 371902 734 372654 856
rect 372822 734 373574 856
rect 373742 734 374494 856
rect 374662 734 375506 856
rect 375674 734 376426 856
rect 376594 734 377346 856
rect 377514 734 378266 856
rect 378434 734 379186 856
rect 379354 734 380106 856
rect 380274 734 381026 856
rect 381194 734 382038 856
rect 382206 734 382958 856
rect 383126 734 383878 856
rect 384046 734 384798 856
rect 384966 734 385718 856
rect 385886 734 386638 856
rect 386806 734 387558 856
rect 387726 734 388570 856
rect 388738 734 389490 856
rect 389658 734 390410 856
rect 390578 734 391330 856
rect 391498 734 392250 856
rect 392418 734 393170 856
rect 393338 734 394090 856
rect 394258 734 395102 856
rect 395270 734 396022 856
rect 396190 734 396942 856
rect 397110 734 397862 856
rect 398030 734 398782 856
rect 398950 734 399702 856
rect 399870 734 400622 856
rect 400790 734 401634 856
rect 401802 734 402554 856
rect 402722 734 403474 856
rect 403642 734 404394 856
rect 404562 734 405314 856
rect 405482 734 406234 856
rect 406402 734 407154 856
rect 407322 734 408166 856
rect 408334 734 409086 856
rect 409254 734 410006 856
rect 410174 734 410926 856
rect 411094 734 411846 856
rect 412014 734 412766 856
rect 412934 734 413686 856
rect 413854 734 414698 856
rect 414866 734 415618 856
rect 415786 734 416538 856
rect 416706 734 417458 856
rect 417626 734 418378 856
rect 418546 734 419298 856
rect 419466 734 420218 856
rect 420386 734 421230 856
rect 421398 734 422150 856
rect 422318 734 423070 856
rect 423238 734 423990 856
rect 424158 734 424910 856
rect 425078 734 425830 856
rect 425998 734 426750 856
rect 426918 734 427762 856
rect 427930 734 428682 856
rect 428850 734 429602 856
rect 429770 734 430522 856
rect 430690 734 431442 856
rect 431610 734 432362 856
rect 432530 734 433282 856
rect 433450 734 434294 856
rect 434462 734 435214 856
rect 435382 734 436134 856
rect 436302 734 437054 856
rect 437222 734 437974 856
rect 438142 734 438894 856
rect 439062 734 439814 856
rect 439982 734 440826 856
rect 440994 734 441746 856
rect 441914 734 442666 856
rect 442834 734 443586 856
rect 443754 734 444506 856
rect 444674 734 445426 856
rect 445594 734 446346 856
rect 446514 734 447358 856
rect 447526 734 448278 856
rect 448446 734 449198 856
rect 449366 734 450118 856
rect 450286 734 451038 856
rect 451206 734 451958 856
rect 452126 734 452878 856
rect 453046 734 453890 856
rect 454058 734 454810 856
rect 454978 734 455730 856
rect 455898 734 456650 856
rect 456818 734 457570 856
rect 457738 734 458490 856
rect 458658 734 459410 856
<< obsm3 >>
rect 4208 2143 449968 457537
<< metal4 >>
rect 4208 2128 4528 457552
rect 19568 2128 19888 457552
rect 34928 2128 35248 457552
rect 50288 2128 50608 457552
rect 65648 2128 65968 457552
rect 81008 2128 81328 457552
rect 96368 2128 96688 457552
rect 111728 2128 112048 457552
rect 127088 2128 127408 457552
rect 142448 2128 142768 457552
rect 157808 2128 158128 457552
rect 173168 2128 173488 457552
rect 188528 2128 188848 457552
rect 203888 2128 204208 457552
rect 219248 2128 219568 457552
rect 234608 2128 234928 457552
rect 249968 2128 250288 457552
rect 265328 2128 265648 457552
rect 280688 2128 281008 457552
rect 296048 2128 296368 457552
rect 311408 2128 311728 457552
rect 326768 2128 327088 457552
rect 342128 2128 342448 457552
rect 357488 2128 357808 457552
rect 372848 2128 373168 457552
rect 388208 2128 388528 457552
rect 403568 2128 403888 457552
rect 418928 2128 419248 457552
rect 434288 2128 434608 457552
rect 449648 2128 449968 457552
<< obsm4 >>
rect 357939 164595 358005 169557
<< labels >>
rlabel metal2 s 1950 459200 2006 460000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 122930 459200 122986 460000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 135074 459200 135130 460000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 147126 459200 147182 460000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 159270 459200 159326 460000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 171414 459200 171470 460000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 183466 459200 183522 460000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 195610 459200 195666 460000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 207662 459200 207718 460000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 219806 459200 219862 460000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 231950 459200 232006 460000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 14002 459200 14058 460000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 244002 459200 244058 460000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 256146 459200 256202 460000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 268198 459200 268254 460000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 280342 459200 280398 460000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 292394 459200 292450 460000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 304538 459200 304594 460000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 316682 459200 316738 460000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 328734 459200 328790 460000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 340878 459200 340934 460000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 352930 459200 352986 460000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 26146 459200 26202 460000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 365074 459200 365130 460000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 377126 459200 377182 460000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 389270 459200 389326 460000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 401414 459200 401470 460000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 413466 459200 413522 460000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 425610 459200 425666 460000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 437662 459200 437718 460000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 449806 459200 449862 460000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 38198 459200 38254 460000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 50342 459200 50398 460000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 62394 459200 62450 460000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 74538 459200 74594 460000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 86682 459200 86738 460000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 98734 459200 98790 460000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 110878 459200 110934 460000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5906 459200 5962 460000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 126978 459200 127034 460000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 139122 459200 139178 460000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 151174 459200 151230 460000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 163318 459200 163374 460000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 175370 459200 175426 460000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 187514 459200 187570 460000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 199658 459200 199714 460000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 211710 459200 211766 460000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 223854 459200 223910 460000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 235906 459200 235962 460000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 18050 459200 18106 460000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 248050 459200 248106 460000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 260194 459200 260250 460000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 272246 459200 272302 460000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 284390 459200 284446 460000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 296442 459200 296498 460000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 308586 459200 308642 460000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 320638 459200 320694 460000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 332782 459200 332838 460000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 344926 459200 344982 460000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 356978 459200 357034 460000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 30194 459200 30250 460000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 369122 459200 369178 460000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 381174 459200 381230 460000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 393318 459200 393374 460000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 405370 459200 405426 460000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 417514 459200 417570 460000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 429658 459200 429714 460000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 441710 459200 441766 460000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 453854 459200 453910 460000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 42246 459200 42302 460000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 54390 459200 54446 460000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 66442 459200 66498 460000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 78586 459200 78642 460000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 90638 459200 90694 460000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 102782 459200 102838 460000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 114926 459200 114982 460000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 9954 459200 10010 460000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 131026 459200 131082 460000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 143170 459200 143226 460000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 155222 459200 155278 460000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 167366 459200 167422 460000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 179418 459200 179474 460000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 191562 459200 191618 460000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 203614 459200 203670 460000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 215758 459200 215814 460000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 227902 459200 227958 460000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 239954 459200 240010 460000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 22098 459200 22154 460000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 252098 459200 252154 460000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 264150 459200 264206 460000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 276294 459200 276350 460000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 288438 459200 288494 460000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 300490 459200 300546 460000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 312634 459200 312690 460000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 324686 459200 324742 460000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 336830 459200 336886 460000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 348882 459200 348938 460000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 361026 459200 361082 460000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 34150 459200 34206 460000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 373170 459200 373226 460000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 385222 459200 385278 460000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 397366 459200 397422 460000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 409418 459200 409474 460000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 421562 459200 421618 460000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 433614 459200 433670 460000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 445758 459200 445814 460000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 457902 459200 457958 460000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 46294 459200 46350 460000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 58438 459200 58494 460000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 70490 459200 70546 460000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 82634 459200 82690 460000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 94686 459200 94742 460000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 106830 459200 106886 460000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 118882 459200 118938 460000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 457626 0 457682 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 458546 0 458602 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 459466 0 459522 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 379242 0 379298 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 382094 0 382150 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 384854 0 384910 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 387614 0 387670 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 390466 0 390522 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 393226 0 393282 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 396078 0 396134 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 398838 0 398894 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 401690 0 401746 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 404450 0 404506 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 407210 0 407266 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 410062 0 410118 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 412822 0 412878 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 415674 0 415730 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 418434 0 418490 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 421286 0 421342 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 424046 0 424102 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 426806 0 426862 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 429658 0 429714 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 432418 0 432474 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 435270 0 435326 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 438030 0 438086 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 440882 0 440938 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 443642 0 443698 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 446402 0 446458 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 449254 0 449310 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 452014 0 452070 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 454866 0 454922 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 174910 0 174966 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 188894 0 188950 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 191746 0 191802 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 197266 0 197322 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 200118 0 200174 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 202878 0 202934 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 205730 0 205786 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 208490 0 208546 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 211342 0 211398 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 214102 0 214158 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 216862 0 216918 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 219714 0 219770 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 225326 0 225382 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 228086 0 228142 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 230938 0 230994 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 233698 0 233754 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 236458 0 236514 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 239310 0 239366 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 242070 0 242126 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 244922 0 244978 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 247682 0 247738 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 253294 0 253350 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 256054 0 256110 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 258906 0 258962 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 261666 0 261722 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 264518 0 264574 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 267278 0 267334 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 270130 0 270186 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 272890 0 272946 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 275650 0 275706 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 278502 0 278558 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 281262 0 281318 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 284114 0 284170 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 286874 0 286930 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 289726 0 289782 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 292486 0 292542 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 295246 0 295302 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 298098 0 298154 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 300858 0 300914 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 303710 0 303766 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 306470 0 306526 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 309230 0 309286 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 312082 0 312138 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 314842 0 314898 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 317694 0 317750 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 320454 0 320510 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 323306 0 323362 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 326066 0 326122 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 328826 0 328882 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 331678 0 331734 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 334438 0 334494 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 337290 0 337346 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 340050 0 340106 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 342902 0 342958 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 345662 0 345718 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 348422 0 348478 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 351274 0 351330 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 354034 0 354090 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 356886 0 356942 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 359646 0 359702 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 362498 0 362554 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 365258 0 365314 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 368018 0 368074 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 370870 0 370926 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 373630 0 373686 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 376482 0 376538 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 380162 0 380218 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 383014 0 383070 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 385774 0 385830 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 388626 0 388682 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 391386 0 391442 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 394146 0 394202 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 396998 0 397054 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 399758 0 399814 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 402610 0 402666 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 405370 0 405426 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 408222 0 408278 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 410982 0 411038 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 413742 0 413798 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 416594 0 416650 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 419354 0 419410 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 422206 0 422262 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 424966 0 425022 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 427818 0 427874 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 430578 0 430634 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 433338 0 433394 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 436190 0 436246 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 438950 0 439006 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 441802 0 441858 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 444562 0 444618 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 447414 0 447470 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 450174 0 450230 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 452934 0 452990 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 455786 0 455842 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 142250 0 142306 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 145102 0 145158 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 147862 0 147918 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 156234 0 156290 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 161846 0 161902 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 164606 0 164662 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 170218 0 170274 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 173070 0 173126 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 178682 0 178738 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 181442 0 181498 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 184202 0 184258 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 187054 0 187110 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 189814 0 189870 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 192666 0 192722 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 195426 0 195482 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 198278 0 198334 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 203798 0 203854 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 206650 0 206706 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 108670 0 108726 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 212262 0 212318 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 215022 0 215078 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 217874 0 217930 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 220634 0 220690 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 223394 0 223450 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 226246 0 226302 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 229006 0 229062 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 231858 0 231914 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 234618 0 234674 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 237470 0 237526 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 240230 0 240286 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 242990 0 243046 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 245842 0 245898 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 248602 0 248658 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 251454 0 251510 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 254214 0 254270 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 257066 0 257122 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 259826 0 259882 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 262586 0 262642 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 265438 0 265494 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 268198 0 268254 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 271050 0 271106 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 273810 0 273866 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 276662 0 276718 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 279422 0 279478 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 282182 0 282238 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 285034 0 285090 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 287794 0 287850 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 290646 0 290702 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 293406 0 293462 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 296258 0 296314 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 299018 0 299074 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 301778 0 301834 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 304630 0 304686 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 307390 0 307446 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 310242 0 310298 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 313002 0 313058 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 315762 0 315818 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 318614 0 318670 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 321374 0 321430 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 324226 0 324282 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 326986 0 327042 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 329838 0 329894 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 332598 0 332654 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 335358 0 335414 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 338210 0 338266 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 340970 0 341026 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 343822 0 343878 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 346582 0 346638 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 349434 0 349490 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 352194 0 352250 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 354954 0 355010 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 357806 0 357862 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 360566 0 360622 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 363418 0 363474 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 366178 0 366234 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 369030 0 369086 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 371790 0 371846 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 374550 0 374606 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 377402 0 377458 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 381082 0 381138 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 383934 0 383990 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 386694 0 386750 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 389546 0 389602 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 392306 0 392362 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 395158 0 395214 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 397918 0 397974 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 400678 0 400734 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 403530 0 403586 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 406290 0 406346 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 409142 0 409198 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 411902 0 411958 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 414754 0 414810 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 417514 0 417570 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 420274 0 420330 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 423126 0 423182 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 425886 0 425942 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 428738 0 428794 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 431498 0 431554 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 434350 0 434406 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 437110 0 437166 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 439870 0 439926 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 442722 0 442778 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 445482 0 445538 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 448334 0 448390 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 451094 0 451150 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 453946 0 454002 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 456706 0 456762 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 182362 0 182418 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 187974 0 188030 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 190734 0 190790 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 193586 0 193642 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 196346 0 196402 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 201958 0 202014 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 207570 0 207626 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 215942 0 215998 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 218794 0 218850 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 224406 0 224462 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 227166 0 227222 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 235538 0 235594 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 238390 0 238446 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 241150 0 241206 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 246762 0 246818 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 249522 0 249578 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 252374 0 252430 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 255134 0 255190 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 257986 0 258042 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 260746 0 260802 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 266358 0 266414 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 269118 0 269174 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 271970 0 272026 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 274730 0 274786 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 280342 0 280398 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 283194 0 283250 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 285954 0 286010 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 288714 0 288770 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 291566 0 291622 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 294326 0 294382 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 297178 0 297234 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 299938 0 299994 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 305550 0 305606 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 308310 0 308366 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 311162 0 311218 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 313922 0 313978 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 316774 0 316830 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 319534 0 319590 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 322294 0 322350 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 325146 0 325202 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 327906 0 327962 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 330758 0 330814 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 333518 0 333574 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 336370 0 336426 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 339130 0 339186 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 341890 0 341946 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 344742 0 344798 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 347502 0 347558 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 350354 0 350410 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 353114 0 353170 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 355966 0 356022 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 358726 0 358782 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 361486 0 361542 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 364338 0 364394 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 367098 0 367154 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 369950 0 370006 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 372710 0 372766 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 375562 0 375618 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 378322 0 378378 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 403568 2128 403888 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 434288 2128 434608 457552 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 418928 2128 419248 457552 6 vssd1
port 503 nsew ground input
rlabel metal4 s 449648 2128 449968 457552 6 vssd1
port 503 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 460000 460000
string LEFview TRUE
string GDS_FILE /project/openlane/computer/runs/computer/results/magic/computer.gds
string GDS_END 102225258
string GDS_START 1009778
<< end >>

