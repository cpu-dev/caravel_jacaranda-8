magic
tech sky130A
magscale 1 2
timestamp 1634795968
<< locali >>
rect 187801 701131 187835 701573
rect 202797 700655 202831 701029
rect 262045 700383 262079 701029
rect 265633 700451 265667 701029
rect 267657 700723 267691 701029
rect 283849 700791 283883 701029
rect 316141 700519 316175 701097
rect 318257 700519 318291 701029
rect 333253 700587 333287 701029
rect 349077 699635 349111 701029
rect 356713 700859 356747 701029
rect 362141 699635 362175 702457
rect 362233 699635 362267 701165
rect 363061 699567 363095 701165
rect 364993 700587 365027 701165
rect 369685 699635 369719 702457
rect 369869 699635 369903 701097
rect 373825 700587 373859 701097
rect 374101 700587 374135 701097
rect 377229 700927 377263 701097
rect 377321 700927 377355 701165
rect 387809 700723 387843 701097
rect 391121 699635 391155 701165
rect 391213 700791 391247 701097
rect 397469 700927 397503 701097
rect 398021 700927 398055 701029
rect 398205 700655 398239 701029
rect 401701 699635 401735 701029
rect 419733 700247 419767 701029
rect 422861 700315 422895 701029
rect 429853 699975 429887 701029
rect 433349 700179 433383 701029
rect 440341 699771 440375 701029
rect 443837 699839 443871 701029
rect 450829 700111 450863 701029
rect 454325 700043 454359 701029
rect 461501 699703 461535 701029
rect 462329 700859 462363 701029
rect 465089 699907 465123 701029
rect 194885 298911 194919 299149
rect 224693 298367 224727 298809
rect 253949 298503 253983 299285
rect 265173 298503 265207 299421
rect 286793 298571 286827 299217
rect 300869 299183 300903 299285
rect 300961 298639 300995 299285
rect 340337 298367 340371 299421
rect 351193 298435 351227 298809
rect 363337 298435 363371 299217
rect 376527 299013 376861 299047
rect 402345 298367 402379 299149
rect 421573 298299 421607 299421
rect 431233 298911 431267 299217
rect 431417 298231 431451 298809
rect 435281 298775 435315 299013
rect 450185 298979 450219 299081
rect 438869 298231 438903 298741
rect 442181 298571 442215 298945
rect 450277 298571 450311 298945
rect 454325 298707 454359 299149
rect 460765 298503 460799 299149
rect 479441 298843 479475 299421
rect 493241 299251 493275 299489
rect 441939 298469 442273 298503
rect 441997 298163 442031 298401
rect 491125 298367 491159 299217
rect 496461 298367 496495 299217
rect 500785 298163 500819 298401
rect 501521 298367 501555 299421
rect 506949 299183 506983 299285
rect 507041 298435 507075 299149
rect 522313 299115 522347 299285
rect 524061 298435 524095 299217
rect 528109 298571 528143 299081
rect 536297 298911 536331 299285
rect 531145 298775 531179 298877
rect 531053 298503 531087 298741
rect 582389 10319 582423 701029
rect 582481 152711 582515 702593
rect 582573 165903 582607 702729
rect 582665 258927 582699 702797
rect 582757 298775 582791 702865
rect 28825 3859 28859 4029
rect 50077 3315 50111 4029
rect 204913 3927 204947 4029
rect 204821 3791 204855 3893
rect 93225 2975 93259 3281
rect 181361 2839 181395 3485
rect 241621 3451 241655 3825
rect 230949 3179 230983 3417
rect 258089 3179 258123 3757
rect 279433 3315 279467 3893
rect 297189 3247 297223 3893
rect 378793 3859 378827 4029
rect 355149 3519 355183 3621
rect 363705 3519 363739 3621
rect 316141 3111 316175 3213
rect 325709 2839 325743 3281
rect 332057 2839 332091 3213
rect 339877 2839 339911 3213
rect 340061 2907 340095 3417
rect 382289 3111 382323 3689
rect 388085 3315 388119 3893
rect 404093 3315 404127 3893
rect 402345 3043 402379 3281
rect 404553 3111 404587 3213
rect 413017 2975 413051 3417
rect 416605 3247 416639 4097
rect 422309 3179 422343 3485
rect 422953 3043 422987 3349
rect 431969 2975 432003 3757
rect 436109 3587 436143 3689
rect 444941 2907 444975 3757
rect 452025 3315 452059 3689
rect 462605 3247 462639 4029
rect 485053 3927 485087 4097
rect 509985 3587 510019 3757
rect 470977 3383 471011 3485
rect 480453 3247 480487 3553
rect 489377 3247 489411 3417
rect 502901 3383 502935 3485
rect 583125 3179 583159 299285
<< viali >>
rect 582757 702865 582791 702899
rect 582665 702797 582699 702831
rect 582573 702729 582607 702763
rect 582481 702593 582515 702627
rect 362141 702457 362175 702491
rect 187801 701573 187835 701607
rect 187801 701097 187835 701131
rect 316141 701097 316175 701131
rect 202797 701029 202831 701063
rect 202797 700621 202831 700655
rect 262045 701029 262079 701063
rect 265633 701029 265667 701063
rect 267657 701029 267691 701063
rect 283849 701029 283883 701063
rect 283849 700757 283883 700791
rect 267657 700689 267691 700723
rect 316141 700485 316175 700519
rect 318257 701029 318291 701063
rect 333253 701029 333287 701063
rect 333253 700553 333287 700587
rect 349077 701029 349111 701063
rect 318257 700485 318291 700519
rect 265633 700417 265667 700451
rect 262045 700349 262079 700383
rect 356713 701029 356747 701063
rect 356713 700825 356747 700859
rect 349077 699601 349111 699635
rect 369685 702457 369719 702491
rect 362141 699601 362175 699635
rect 362233 701165 362267 701199
rect 362233 699601 362267 699635
rect 363061 701165 363095 701199
rect 364993 701165 365027 701199
rect 364993 700553 365027 700587
rect 377321 701165 377355 701199
rect 369685 699601 369719 699635
rect 369869 701097 369903 701131
rect 373825 701097 373859 701131
rect 373825 700553 373859 700587
rect 374101 701097 374135 701131
rect 377229 701097 377263 701131
rect 377229 700893 377263 700927
rect 391121 701165 391155 701199
rect 377321 700893 377355 700927
rect 387809 701097 387843 701131
rect 387809 700689 387843 700723
rect 374101 700553 374135 700587
rect 369869 699601 369903 699635
rect 391213 701097 391247 701131
rect 397469 701097 397503 701131
rect 397469 700893 397503 700927
rect 398021 701029 398055 701063
rect 398021 700893 398055 700927
rect 398205 701029 398239 701063
rect 391213 700757 391247 700791
rect 398205 700621 398239 700655
rect 401701 701029 401735 701063
rect 391121 699601 391155 699635
rect 419733 701029 419767 701063
rect 422861 701029 422895 701063
rect 422861 700281 422895 700315
rect 429853 701029 429887 701063
rect 419733 700213 419767 700247
rect 433349 701029 433383 701063
rect 433349 700145 433383 700179
rect 440341 701029 440375 701063
rect 429853 699941 429887 699975
rect 443837 701029 443871 701063
rect 450829 701029 450863 701063
rect 450829 700077 450863 700111
rect 454325 701029 454359 701063
rect 454325 700009 454359 700043
rect 461501 701029 461535 701063
rect 443837 699805 443871 699839
rect 440341 699737 440375 699771
rect 462329 701029 462363 701063
rect 462329 700825 462363 700859
rect 465089 701029 465123 701063
rect 465089 699873 465123 699907
rect 582389 701029 582423 701063
rect 461501 699669 461535 699703
rect 401701 699601 401735 699635
rect 363061 699533 363095 699567
rect 493241 299489 493275 299523
rect 265173 299421 265207 299455
rect 253949 299285 253983 299319
rect 194885 299149 194919 299183
rect 194885 298877 194919 298911
rect 224693 298809 224727 298843
rect 253949 298469 253983 298503
rect 340337 299421 340371 299455
rect 300869 299285 300903 299319
rect 286793 299217 286827 299251
rect 300869 299149 300903 299183
rect 300961 299285 300995 299319
rect 300961 298605 300995 298639
rect 286793 298537 286827 298571
rect 265173 298469 265207 298503
rect 224693 298333 224727 298367
rect 421573 299421 421607 299455
rect 363337 299217 363371 299251
rect 351193 298809 351227 298843
rect 351193 298401 351227 298435
rect 402345 299149 402379 299183
rect 376493 299013 376527 299047
rect 376861 299013 376895 299047
rect 363337 298401 363371 298435
rect 340337 298333 340371 298367
rect 402345 298333 402379 298367
rect 479441 299421 479475 299455
rect 431233 299217 431267 299251
rect 454325 299149 454359 299183
rect 450185 299081 450219 299115
rect 431233 298877 431267 298911
rect 435281 299013 435315 299047
rect 421573 298265 421607 298299
rect 431417 298809 431451 298843
rect 442181 298945 442215 298979
rect 450185 298945 450219 298979
rect 450277 298945 450311 298979
rect 435281 298741 435315 298775
rect 438869 298741 438903 298775
rect 431417 298197 431451 298231
rect 442181 298537 442215 298571
rect 454325 298673 454359 298707
rect 460765 299149 460799 299183
rect 450277 298537 450311 298571
rect 501521 299421 501555 299455
rect 479441 298809 479475 298843
rect 491125 299217 491159 299251
rect 493241 299217 493275 299251
rect 496461 299217 496495 299251
rect 441905 298469 441939 298503
rect 442273 298469 442307 298503
rect 460765 298469 460799 298503
rect 438869 298197 438903 298231
rect 441997 298401 442031 298435
rect 491125 298333 491159 298367
rect 496461 298333 496495 298367
rect 500785 298401 500819 298435
rect 441997 298129 442031 298163
rect 506949 299285 506983 299319
rect 522313 299285 522347 299319
rect 506949 299149 506983 299183
rect 507041 299149 507075 299183
rect 536297 299285 536331 299319
rect 522313 299081 522347 299115
rect 524061 299217 524095 299251
rect 507041 298401 507075 298435
rect 528109 299081 528143 299115
rect 531145 298877 531179 298911
rect 536297 298877 536331 298911
rect 528109 298537 528143 298571
rect 531053 298741 531087 298775
rect 531145 298741 531179 298775
rect 531053 298469 531087 298503
rect 524061 298401 524095 298435
rect 501521 298333 501555 298367
rect 500785 298129 500819 298163
rect 582757 298741 582791 298775
rect 583125 299285 583159 299319
rect 582665 258893 582699 258927
rect 582573 165869 582607 165903
rect 582481 152677 582515 152711
rect 582389 10285 582423 10319
rect 416605 4097 416639 4131
rect 28825 4029 28859 4063
rect 28825 3825 28859 3859
rect 50077 4029 50111 4063
rect 204913 4029 204947 4063
rect 378793 4029 378827 4063
rect 204821 3893 204855 3927
rect 204913 3893 204947 3927
rect 279433 3893 279467 3927
rect 204821 3757 204855 3791
rect 241621 3825 241655 3859
rect 181361 3485 181395 3519
rect 50077 3281 50111 3315
rect 93225 3281 93259 3315
rect 93225 2941 93259 2975
rect 230949 3417 230983 3451
rect 241621 3417 241655 3451
rect 258089 3757 258123 3791
rect 230949 3145 230983 3179
rect 279433 3281 279467 3315
rect 297189 3893 297223 3927
rect 378793 3825 378827 3859
rect 388085 3893 388119 3927
rect 382289 3689 382323 3723
rect 355149 3621 355183 3655
rect 355149 3485 355183 3519
rect 363705 3621 363739 3655
rect 363705 3485 363739 3519
rect 340061 3417 340095 3451
rect 325709 3281 325743 3315
rect 297189 3213 297223 3247
rect 316141 3213 316175 3247
rect 258089 3145 258123 3179
rect 316141 3077 316175 3111
rect 181361 2805 181395 2839
rect 325709 2805 325743 2839
rect 332057 3213 332091 3247
rect 332057 2805 332091 2839
rect 339877 3213 339911 3247
rect 404093 3893 404127 3927
rect 388085 3281 388119 3315
rect 402345 3281 402379 3315
rect 404093 3281 404127 3315
rect 413017 3417 413051 3451
rect 382289 3077 382323 3111
rect 404553 3213 404587 3247
rect 404553 3077 404587 3111
rect 402345 3009 402379 3043
rect 485053 4097 485087 4131
rect 462605 4029 462639 4063
rect 431969 3757 432003 3791
rect 416605 3213 416639 3247
rect 422309 3485 422343 3519
rect 422309 3145 422343 3179
rect 422953 3349 422987 3383
rect 422953 3009 422987 3043
rect 413017 2941 413051 2975
rect 444941 3757 444975 3791
rect 436109 3689 436143 3723
rect 436109 3553 436143 3587
rect 431969 2941 432003 2975
rect 340061 2873 340095 2907
rect 452025 3689 452059 3723
rect 452025 3281 452059 3315
rect 485053 3893 485087 3927
rect 509985 3757 510019 3791
rect 480453 3553 480487 3587
rect 509985 3553 510019 3587
rect 470977 3485 471011 3519
rect 470977 3349 471011 3383
rect 462605 3213 462639 3247
rect 502901 3485 502935 3519
rect 480453 3213 480487 3247
rect 489377 3417 489411 3451
rect 502901 3349 502935 3383
rect 489377 3213 489411 3247
rect 583125 3145 583159 3179
rect 444941 2873 444975 2907
rect 339877 2805 339911 2839
<< metal1 >>
rect 15838 703740 15844 703792
rect 15896 703780 15902 703792
rect 552934 703780 552940 703792
rect 15896 703752 552940 703780
rect 15896 703740 15902 703752
rect 552934 703740 552940 703752
rect 552992 703740 552998 703792
rect 22738 703672 22744 703724
rect 22796 703712 22802 703724
rect 563514 703712 563520 703724
rect 22796 703684 563520 703712
rect 22796 703672 22802 703684
rect 563514 703672 563520 703684
rect 563572 703672 563578 703724
rect 363506 703604 363512 703656
rect 363564 703644 363570 703656
rect 429654 703644 429660 703656
rect 363564 703616 429660 703644
rect 363564 703604 363570 703616
rect 429654 703604 429660 703616
rect 429712 703604 429718 703656
rect 300302 703536 300308 703588
rect 300360 703576 300366 703588
rect 384574 703576 384580 703588
rect 300360 703548 384580 703576
rect 300360 703536 300366 703548
rect 384574 703536 384580 703548
rect 384632 703536 384638 703588
rect 374546 703468 374552 703520
rect 374604 703508 374610 703520
rect 577038 703508 577044 703520
rect 374604 703480 577044 703508
rect 374604 703468 374610 703480
rect 577038 703468 577044 703480
rect 577096 703468 577102 703520
rect 182174 703400 182180 703452
rect 182232 703440 182238 703452
rect 437198 703440 437204 703452
rect 182232 703412 437204 703440
rect 182232 703400 182238 703412
rect 437198 703400 437204 703412
rect 437256 703400 437262 703452
rect 349430 703332 349436 703384
rect 349488 703372 349494 703384
rect 543458 703372 543464 703384
rect 349488 703344 543464 703372
rect 349488 703332 349494 703344
rect 543458 703332 543464 703344
rect 543516 703332 543522 703384
rect 182266 703264 182272 703316
rect 182324 703304 182330 703316
rect 447686 703304 447692 703316
rect 182324 703276 447692 703304
rect 182324 703264 182330 703276
rect 447686 703264 447692 703276
rect 447744 703264 447750 703316
rect 182358 703196 182364 703248
rect 182416 703236 182422 703248
rect 458174 703236 458180 703248
rect 182416 703208 458180 703236
rect 182416 703196 182422 703208
rect 458174 703196 458180 703208
rect 458232 703196 458238 703248
rect 182450 703128 182456 703180
rect 182508 703168 182514 703180
rect 468754 703168 468760 703180
rect 182508 703140 468760 703168
rect 182508 703128 182514 703140
rect 468754 703128 468760 703140
rect 468812 703128 468818 703180
rect 182542 703060 182548 703112
rect 182600 703100 182606 703112
rect 479242 703100 479248 703112
rect 182600 703072 479248 703100
rect 182600 703060 182606 703072
rect 479242 703060 479248 703072
rect 479300 703060 479306 703112
rect 182634 702992 182640 703044
rect 182692 703032 182698 703044
rect 489822 703032 489828 703044
rect 182692 703004 489828 703032
rect 182692 702992 182698 703004
rect 489822 702992 489828 703004
rect 489880 702992 489886 703044
rect 182726 702924 182732 702976
rect 182784 702964 182790 702976
rect 500310 702964 500316 702976
rect 182784 702936 500316 702964
rect 182784 702924 182790 702936
rect 500310 702924 500316 702936
rect 500368 702924 500374 702976
rect 258166 702856 258172 702908
rect 258224 702896 258230 702908
rect 582745 702899 582803 702905
rect 582745 702896 582757 702899
rect 258224 702868 582757 702896
rect 258224 702856 258230 702868
rect 582745 702865 582757 702868
rect 582791 702865 582803 702899
rect 582745 702859 582803 702865
rect 254670 702788 254676 702840
rect 254728 702828 254734 702840
rect 582653 702831 582711 702837
rect 582653 702828 582665 702831
rect 254728 702800 582665 702828
rect 254728 702788 254734 702800
rect 582653 702797 582665 702800
rect 582699 702797 582711 702831
rect 582653 702791 582711 702797
rect 226610 702720 226616 702772
rect 226668 702760 226674 702772
rect 582561 702763 582619 702769
rect 582561 702760 582573 702763
rect 226668 702732 582573 702760
rect 226668 702720 226674 702732
rect 582561 702729 582573 702732
rect 582607 702729 582619 702763
rect 582561 702723 582619 702729
rect 180058 702652 180064 702704
rect 180116 702692 180122 702704
rect 542446 702692 542452 702704
rect 180116 702664 542452 702692
rect 180116 702652 180122 702664
rect 542446 702652 542452 702664
rect 542504 702652 542510 702704
rect 219618 702584 219624 702636
rect 219676 702624 219682 702636
rect 582469 702627 582527 702633
rect 582469 702624 582481 702627
rect 219676 702596 582481 702624
rect 219676 702584 219682 702596
rect 582469 702593 582481 702596
rect 582515 702593 582527 702627
rect 582469 702587 582527 702593
rect 300302 702516 300308 702568
rect 300360 702556 300366 702568
rect 375374 702556 375380 702568
rect 300360 702528 375380 702556
rect 300360 702516 300366 702528
rect 375374 702516 375380 702528
rect 375432 702516 375438 702568
rect 404354 702516 404360 702568
rect 404412 702556 404418 702568
rect 409046 702556 409052 702568
rect 404412 702528 409052 702556
rect 404412 702516 404418 702528
rect 409046 702516 409052 702528
rect 409104 702516 409110 702568
rect 362129 702491 362187 702497
rect 362129 702457 362141 702491
rect 362175 702488 362187 702491
rect 365714 702488 365720 702500
rect 362175 702460 365720 702488
rect 362175 702457 362187 702460
rect 362129 702451 362187 702457
rect 365714 702448 365720 702460
rect 365772 702448 365778 702500
rect 369670 702488 369676 702500
rect 369631 702460 369676 702488
rect 369670 702448 369676 702460
rect 369728 702448 369734 702500
rect 370498 702448 370504 702500
rect 370556 702488 370562 702500
rect 413646 702488 413652 702500
rect 370556 702460 413652 702488
rect 370556 702448 370562 702460
rect 413646 702448 413652 702460
rect 413704 702448 413710 702500
rect 35158 702380 35164 702432
rect 35216 702420 35222 702432
rect 486326 702420 486332 702432
rect 35216 702392 486332 702420
rect 35216 702380 35222 702392
rect 486326 702380 486332 702392
rect 486384 702380 486390 702432
rect 18598 702312 18604 702364
rect 18656 702352 18662 702364
rect 475746 702352 475752 702364
rect 18656 702324 475752 702352
rect 18656 702312 18662 702324
rect 475746 702312 475752 702324
rect 475804 702312 475810 702364
rect 14458 702244 14464 702296
rect 14516 702284 14522 702296
rect 472250 702284 472256 702296
rect 14516 702256 472256 702284
rect 14516 702244 14522 702256
rect 472250 702244 472256 702256
rect 472308 702244 472314 702296
rect 289814 702176 289820 702228
rect 289872 702216 289878 702228
rect 333974 702216 333980 702228
rect 289872 702188 333980 702216
rect 289872 702176 289878 702188
rect 333974 702176 333980 702188
rect 334032 702176 334038 702228
rect 338942 702176 338948 702228
rect 339000 702216 339006 702228
rect 427630 702216 427636 702228
rect 339000 702188 427636 702216
rect 339000 702176 339006 702188
rect 427630 702176 427636 702188
rect 427688 702176 427694 702228
rect 314378 702108 314384 702160
rect 314436 702148 314442 702160
rect 418062 702148 418068 702160
rect 314436 702120 418068 702148
rect 314436 702108 314442 702120
rect 418062 702108 418068 702120
rect 418120 702108 418126 702160
rect 268746 702040 268752 702092
rect 268804 702080 268810 702092
rect 374546 702080 374552 702092
rect 268804 702052 374552 702080
rect 268804 702040 268810 702052
rect 374546 702040 374552 702052
rect 374604 702040 374610 702092
rect 374638 702040 374644 702092
rect 374696 702080 374702 702092
rect 556430 702080 556436 702092
rect 374696 702052 556436 702080
rect 374696 702040 374702 702052
rect 556430 702040 556436 702052
rect 556488 702040 556494 702092
rect 328362 701972 328368 702024
rect 328420 702012 328426 702024
rect 583754 702012 583760 702024
rect 328420 701984 583760 702012
rect 328420 701972 328426 701984
rect 583754 701972 583760 701984
rect 583812 701972 583818 702024
rect 324866 701904 324872 701956
rect 324924 701944 324930 701956
rect 583846 701944 583852 701956
rect 324924 701916 583852 701944
rect 324924 701904 324930 701916
rect 583846 701904 583852 701916
rect 583904 701904 583910 701956
rect 307294 701836 307300 701888
rect 307352 701876 307358 701888
rect 583570 701876 583576 701888
rect 307352 701848 583576 701876
rect 307352 701836 307358 701848
rect 583570 701836 583576 701848
rect 583628 701836 583634 701888
rect 304074 701768 304080 701820
rect 304132 701808 304138 701820
rect 582558 701808 582564 701820
rect 304132 701780 582564 701808
rect 304132 701768 304138 701780
rect 582558 701768 582564 701780
rect 582616 701768 582622 701820
rect 181806 701700 181812 701752
rect 181864 701740 181870 701752
rect 181864 701712 190454 701740
rect 181864 701700 181870 701712
rect 182082 701632 182088 701684
rect 182140 701672 182146 701684
rect 190426 701672 190454 701712
rect 297082 701700 297088 701752
rect 297140 701740 297146 701752
rect 583386 701740 583392 701752
rect 297140 701712 583392 701740
rect 297140 701700 297146 701712
rect 583386 701700 583392 701712
rect 583444 701700 583450 701752
rect 201678 701672 201684 701684
rect 182140 701644 187924 701672
rect 190426 701644 201684 701672
rect 182140 701632 182146 701644
rect 181898 701564 181904 701616
rect 181956 701604 181962 701616
rect 187789 701607 187847 701613
rect 187789 701604 187801 701607
rect 181956 701576 187801 701604
rect 181956 701564 181962 701576
rect 187789 701573 187801 701576
rect 187835 701573 187847 701607
rect 187896 701604 187924 701644
rect 201678 701632 201684 701644
rect 201736 701632 201742 701684
rect 293586 701632 293592 701684
rect 293644 701672 293650 701684
rect 583478 701672 583484 701684
rect 293644 701644 583484 701672
rect 293644 701632 293650 701644
rect 583478 701632 583484 701644
rect 583536 701632 583542 701684
rect 191190 701604 191196 701616
rect 187896 701576 191196 701604
rect 187789 701567 187847 701573
rect 191190 701564 191196 701576
rect 191248 701564 191254 701616
rect 286594 701564 286600 701616
rect 286652 701604 286658 701616
rect 583202 701604 583208 701616
rect 286652 701576 583208 701604
rect 286652 701564 286658 701576
rect 583202 701564 583208 701576
rect 583260 701564 583266 701616
rect 183002 701496 183008 701548
rect 183060 701536 183066 701548
rect 205174 701536 205180 701548
rect 183060 701508 205180 701536
rect 183060 701496 183066 701508
rect 205174 701496 205180 701508
rect 205232 701496 205238 701548
rect 282822 701496 282828 701548
rect 282880 701536 282886 701548
rect 583294 701536 583300 701548
rect 282880 701508 583300 701536
rect 282880 701496 282886 701508
rect 583294 701496 583300 701508
rect 583352 701496 583358 701548
rect 182910 701428 182916 701480
rect 182968 701468 182974 701480
rect 208670 701468 208676 701480
rect 182968 701440 208676 701468
rect 182968 701428 182974 701440
rect 208670 701428 208676 701440
rect 208728 701428 208734 701480
rect 279602 701428 279608 701480
rect 279660 701468 279666 701480
rect 583110 701468 583116 701480
rect 279660 701440 583116 701468
rect 279660 701428 279666 701440
rect 583110 701428 583116 701440
rect 583168 701428 583174 701480
rect 137278 701360 137284 701412
rect 137336 701400 137342 701412
rect 243998 701400 244004 701412
rect 137336 701372 244004 701400
rect 137336 701360 137342 701372
rect 243998 701360 244004 701372
rect 244056 701360 244062 701412
rect 275922 701360 275928 701412
rect 275980 701400 275986 701412
rect 582926 701400 582932 701412
rect 275980 701372 582932 701400
rect 275980 701360 275986 701372
rect 582926 701360 582932 701372
rect 582984 701360 582990 701412
rect 39298 701292 39304 701344
rect 39356 701332 39362 701344
rect 247862 701332 247868 701344
rect 39356 701304 247868 701332
rect 39356 701292 39362 701304
rect 247862 701292 247868 701304
rect 247920 701292 247926 701344
rect 272610 701292 272616 701344
rect 272668 701332 272674 701344
rect 583018 701332 583024 701344
rect 272668 701304 583024 701332
rect 272668 701292 272674 701304
rect 583018 701292 583024 701304
rect 583076 701292 583082 701344
rect 32398 701224 32404 701276
rect 32456 701264 32462 701276
rect 482462 701264 482468 701276
rect 32456 701236 482468 701264
rect 32456 701224 32462 701236
rect 482462 701224 482468 701236
rect 482520 701224 482526 701276
rect 183094 701156 183100 701208
rect 183152 701196 183158 701208
rect 194686 701196 194692 701208
rect 183152 701168 194692 701196
rect 183152 701156 183158 701168
rect 194686 701156 194692 701168
rect 194744 701156 194750 701208
rect 362218 701196 362224 701208
rect 362179 701168 362224 701196
rect 362218 701156 362224 701168
rect 362276 701156 362282 701208
rect 362954 701156 362960 701208
rect 363012 701196 363018 701208
rect 363049 701199 363107 701205
rect 363049 701196 363061 701199
rect 363012 701168 363061 701196
rect 363012 701156 363018 701168
rect 363049 701165 363061 701168
rect 363095 701165 363107 701199
rect 364978 701196 364984 701208
rect 364939 701168 364984 701196
rect 363049 701159 363107 701165
rect 364978 701156 364984 701168
rect 365036 701156 365042 701208
rect 367094 701156 367100 701208
rect 367152 701196 367158 701208
rect 377309 701199 377367 701205
rect 377309 701196 377321 701199
rect 367152 701168 377321 701196
rect 367152 701156 367158 701168
rect 377309 701165 377321 701168
rect 377355 701165 377367 701199
rect 391106 701196 391112 701208
rect 391067 701168 391112 701196
rect 377309 701159 377367 701165
rect 391106 701156 391112 701168
rect 391164 701156 391170 701208
rect 532234 701156 532240 701208
rect 532292 701196 532298 701208
rect 535546 701196 535552 701208
rect 532292 701168 535552 701196
rect 532292 701156 532298 701168
rect 535546 701156 535552 701168
rect 535604 701156 535610 701208
rect 181990 701088 181996 701140
rect 182048 701128 182054 701140
rect 187694 701128 187700 701140
rect 182048 701100 187700 701128
rect 182048 701088 182054 701100
rect 187694 701088 187700 701100
rect 187752 701088 187758 701140
rect 187789 701131 187847 701137
rect 187789 701097 187801 701131
rect 187835 701128 187847 701131
rect 198182 701128 198188 701140
rect 187835 701100 198188 701128
rect 187835 701097 187847 701100
rect 187789 701091 187847 701097
rect 198182 701088 198188 701100
rect 198240 701088 198246 701140
rect 316126 701128 316132 701140
rect 316087 701100 316132 701128
rect 316126 701088 316132 701100
rect 316184 701088 316190 701140
rect 332428 701100 332640 701128
rect 182818 701020 182824 701072
rect 182876 701060 182882 701072
rect 184198 701060 184204 701072
rect 182876 701032 184204 701060
rect 182876 701020 182882 701032
rect 184198 701020 184204 701032
rect 184256 701020 184262 701072
rect 202782 701060 202788 701072
rect 202743 701032 202788 701060
rect 202782 701020 202788 701032
rect 202840 701020 202846 701072
rect 262030 701060 262036 701072
rect 261991 701032 262036 701060
rect 262030 701020 262036 701032
rect 262088 701020 262094 701072
rect 265618 701060 265624 701072
rect 265579 701032 265624 701060
rect 265618 701020 265624 701032
rect 265676 701020 265682 701072
rect 267642 701060 267648 701072
rect 267603 701032 267648 701060
rect 267642 701020 267648 701032
rect 267700 701020 267706 701072
rect 283834 701060 283840 701072
rect 283795 701032 283840 701060
rect 283834 701020 283840 701032
rect 283892 701020 283898 701072
rect 318242 701060 318248 701072
rect 318203 701032 318248 701060
rect 318242 701020 318248 701032
rect 318300 701020 318306 701072
rect 137830 700952 137836 701004
rect 137888 700992 137894 701004
rect 332428 700992 332456 701100
rect 332502 701020 332508 701072
rect 332560 701020 332566 701072
rect 137888 700964 332456 700992
rect 137888 700952 137894 700964
rect 332520 700924 332548 701020
rect 332612 700992 332640 701100
rect 335722 701088 335728 701140
rect 335780 701128 335786 701140
rect 365806 701128 365812 701140
rect 335780 701100 365812 701128
rect 335780 701088 335786 701100
rect 365806 701088 365812 701100
rect 365864 701088 365870 701140
rect 369486 701088 369492 701140
rect 369544 701128 369550 701140
rect 369857 701131 369915 701137
rect 369857 701128 369869 701131
rect 369544 701100 369869 701128
rect 369544 701088 369550 701100
rect 369857 701097 369869 701100
rect 369903 701097 369915 701131
rect 373810 701128 373816 701140
rect 373771 701100 373816 701128
rect 369857 701091 369915 701097
rect 373810 701088 373816 701100
rect 373868 701088 373874 701140
rect 374086 701128 374092 701140
rect 374047 701100 374092 701128
rect 374086 701088 374092 701100
rect 374144 701088 374150 701140
rect 377214 701128 377220 701140
rect 377175 701100 377220 701128
rect 377214 701088 377220 701100
rect 377272 701088 377278 701140
rect 387794 701128 387800 701140
rect 387755 701100 387800 701128
rect 387794 701088 387800 701100
rect 387852 701088 387858 701140
rect 391198 701128 391204 701140
rect 391159 701100 391204 701128
rect 391198 701088 391204 701100
rect 391256 701088 391262 701140
rect 397454 701128 397460 701140
rect 397415 701100 397460 701128
rect 397454 701088 397460 701100
rect 397512 701088 397518 701140
rect 333238 701060 333244 701072
rect 333199 701032 333244 701060
rect 333238 701020 333244 701032
rect 333296 701020 333302 701072
rect 349062 701060 349068 701072
rect 349023 701032 349068 701060
rect 349062 701020 349068 701032
rect 349120 701020 349126 701072
rect 356698 701060 356704 701072
rect 356659 701032 356704 701060
rect 356698 701020 356704 701032
rect 356756 701020 356762 701072
rect 360102 701020 360108 701072
rect 360160 701060 360166 701072
rect 398009 701063 398067 701069
rect 398009 701060 398021 701063
rect 360160 701032 398021 701060
rect 360160 701020 360166 701032
rect 398009 701029 398021 701032
rect 398055 701029 398067 701063
rect 398190 701060 398196 701072
rect 398151 701032 398196 701060
rect 398009 701023 398067 701029
rect 398190 701020 398196 701032
rect 398248 701020 398254 701072
rect 401686 701060 401692 701072
rect 401647 701032 401692 701060
rect 401686 701020 401692 701032
rect 401744 701020 401750 701072
rect 404354 701020 404360 701072
rect 404412 701020 404418 701072
rect 419718 701060 419724 701072
rect 419679 701032 419724 701060
rect 419718 701020 419724 701032
rect 419776 701020 419782 701072
rect 422846 701060 422852 701072
rect 422807 701032 422852 701060
rect 422846 701020 422852 701032
rect 422904 701020 422910 701072
rect 429838 701060 429844 701072
rect 429799 701032 429844 701060
rect 429838 701020 429844 701032
rect 429896 701020 429902 701072
rect 433334 701060 433340 701072
rect 433295 701032 433340 701060
rect 433334 701020 433340 701032
rect 433392 701020 433398 701072
rect 440326 701060 440332 701072
rect 440287 701032 440332 701060
rect 440326 701020 440332 701032
rect 440384 701020 440390 701072
rect 443822 701060 443828 701072
rect 443783 701032 443828 701060
rect 443822 701020 443828 701032
rect 443880 701020 443886 701072
rect 450814 701060 450820 701072
rect 450775 701032 450820 701060
rect 450814 701020 450820 701032
rect 450872 701020 450878 701072
rect 454310 701060 454316 701072
rect 454271 701032 454316 701060
rect 454310 701020 454316 701032
rect 454368 701020 454374 701072
rect 461486 701060 461492 701072
rect 461447 701032 461492 701060
rect 461486 701020 461492 701032
rect 461544 701020 461550 701072
rect 462314 701060 462320 701072
rect 462275 701032 462320 701060
rect 462314 701020 462320 701032
rect 462372 701020 462378 701072
rect 465074 701060 465080 701072
rect 465035 701032 465080 701060
rect 465074 701020 465080 701032
rect 465132 701020 465138 701072
rect 478506 701020 478512 701072
rect 478564 701020 478570 701072
rect 566734 701020 566740 701072
rect 566792 701020 566798 701072
rect 577866 701020 577872 701072
rect 577924 701060 577930 701072
rect 582377 701063 582435 701069
rect 582377 701060 582389 701063
rect 577924 701032 582389 701060
rect 577924 701020 577930 701032
rect 582377 701029 582389 701032
rect 582423 701029 582435 701063
rect 582377 701023 582435 701029
rect 404372 700992 404400 701020
rect 332612 700964 404400 700992
rect 377217 700927 377275 700933
rect 377217 700924 377229 700927
rect 332520 700896 377229 700924
rect 377217 700893 377229 700896
rect 377263 700893 377275 700927
rect 377217 700887 377275 700893
rect 377309 700927 377367 700933
rect 377309 700893 377321 700927
rect 377355 700924 377367 700927
rect 397457 700927 397515 700933
rect 397457 700924 397469 700927
rect 377355 700896 397469 700924
rect 377355 700893 377367 700896
rect 377309 700887 377367 700893
rect 397457 700893 397469 700896
rect 397503 700893 397515 700927
rect 397457 700887 397515 700893
rect 398009 700927 398067 700933
rect 398009 700893 398021 700927
rect 398055 700924 398067 700927
rect 478524 700924 478552 701020
rect 398055 700896 478552 700924
rect 398055 700893 398067 700896
rect 398009 700887 398067 700893
rect 356701 700859 356759 700865
rect 356701 700825 356713 700859
rect 356747 700856 356759 700859
rect 462317 700859 462375 700865
rect 462317 700856 462329 700859
rect 356747 700828 462329 700856
rect 356747 700825 356759 700828
rect 356701 700819 356759 700825
rect 462317 700825 462329 700828
rect 462363 700825 462375 700859
rect 462317 700819 462375 700825
rect 283837 700791 283895 700797
rect 283837 700757 283849 700791
rect 283883 700788 283895 700791
rect 391201 700791 391259 700797
rect 391201 700788 391213 700791
rect 283883 700760 391213 700788
rect 283883 700757 283895 700760
rect 283837 700751 283895 700757
rect 391201 700757 391213 700760
rect 391247 700757 391259 700791
rect 391201 700751 391259 700757
rect 267645 700723 267703 700729
rect 267645 700689 267657 700723
rect 267691 700720 267703 700723
rect 387797 700723 387855 700729
rect 387797 700720 387809 700723
rect 267691 700692 387809 700720
rect 267691 700689 267703 700692
rect 267645 700683 267703 700689
rect 387797 700689 387809 700692
rect 387843 700689 387855 700723
rect 387797 700683 387855 700689
rect 202785 700655 202843 700661
rect 202785 700621 202797 700655
rect 202831 700652 202843 700655
rect 398193 700655 398251 700661
rect 398193 700652 398205 700655
rect 202831 700624 398205 700652
rect 202831 700621 202843 700624
rect 202785 700615 202843 700621
rect 398193 700621 398205 700624
rect 398239 700621 398251 700655
rect 398193 700615 398251 700621
rect 61378 700544 61384 700596
rect 61436 700584 61442 700596
rect 333241 700587 333299 700593
rect 333241 700584 333253 700587
rect 61436 700556 333253 700584
rect 61436 700544 61442 700556
rect 333241 700553 333253 700556
rect 333287 700553 333299 700587
rect 333241 700547 333299 700553
rect 364981 700587 365039 700593
rect 364981 700553 364993 700587
rect 365027 700584 365039 700587
rect 373813 700587 373871 700593
rect 373813 700584 373825 700587
rect 365027 700556 373825 700584
rect 365027 700553 365039 700556
rect 364981 700547 365039 700553
rect 373813 700553 373825 700556
rect 373859 700553 373871 700587
rect 373813 700547 373871 700553
rect 374089 700587 374147 700593
rect 374089 700553 374101 700587
rect 374135 700584 374147 700587
rect 566752 700584 566780 701020
rect 374135 700556 566780 700584
rect 374135 700553 374147 700556
rect 374089 700547 374147 700553
rect 36538 700476 36544 700528
rect 36596 700516 36602 700528
rect 316129 700519 316187 700525
rect 316129 700516 316141 700519
rect 36596 700488 316141 700516
rect 36596 700476 36602 700488
rect 316129 700485 316141 700488
rect 316175 700485 316187 700519
rect 316129 700479 316187 700485
rect 318245 700519 318303 700525
rect 318245 700485 318257 700519
rect 318291 700516 318303 700519
rect 583662 700516 583668 700528
rect 318291 700488 583668 700516
rect 318291 700485 318303 700488
rect 318245 700479 318303 700485
rect 583662 700476 583668 700488
rect 583720 700476 583726 700528
rect 265621 700451 265679 700457
rect 265621 700417 265633 700451
rect 265667 700448 265679 700451
rect 582742 700448 582748 700460
rect 265667 700420 582748 700448
rect 265667 700417 265679 700420
rect 265621 700411 265679 700417
rect 582742 700408 582748 700420
rect 582800 700408 582806 700460
rect 262033 700383 262091 700389
rect 262033 700349 262045 700383
rect 262079 700380 262091 700383
rect 582834 700380 582840 700392
rect 262079 700352 582840 700380
rect 262079 700349 262091 700352
rect 262033 700343 262091 700349
rect 582834 700340 582840 700352
rect 582892 700340 582898 700392
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 422849 700315 422907 700321
rect 422849 700312 422861 700315
rect 89220 700284 422861 700312
rect 89220 700272 89226 700284
rect 422849 700281 422861 700284
rect 422895 700281 422907 700315
rect 422849 700275 422907 700281
rect 72970 700204 72976 700256
rect 73028 700244 73034 700256
rect 419721 700247 419779 700253
rect 419721 700244 419733 700247
rect 73028 700216 419733 700244
rect 73028 700204 73034 700216
rect 419721 700213 419733 700216
rect 419767 700213 419779 700247
rect 419721 700207 419779 700213
rect 24302 700136 24308 700188
rect 24360 700176 24366 700188
rect 433337 700179 433395 700185
rect 433337 700176 433349 700179
rect 24360 700148 433349 700176
rect 24360 700136 24366 700148
rect 433337 700145 433349 700148
rect 433383 700145 433395 700179
rect 433337 700139 433395 700145
rect 32490 700068 32496 700120
rect 32548 700108 32554 700120
rect 450817 700111 450875 700117
rect 450817 700108 450829 700111
rect 32548 700080 450829 700108
rect 32548 700068 32554 700080
rect 450817 700077 450829 700080
rect 450863 700077 450875 700111
rect 450817 700071 450875 700077
rect 35250 700000 35256 700052
rect 35308 700040 35314 700052
rect 454313 700043 454371 700049
rect 454313 700040 454325 700043
rect 35308 700012 454325 700040
rect 35308 700000 35314 700012
rect 454313 700009 454325 700012
rect 454359 700009 454371 700043
rect 454313 700003 454371 700009
rect 8110 699932 8116 699984
rect 8168 699972 8174 699984
rect 429841 699975 429899 699981
rect 429841 699972 429853 699975
rect 8168 699944 429853 699972
rect 8168 699932 8174 699944
rect 429841 699941 429853 699944
rect 429887 699941 429899 699975
rect 429841 699935 429899 699941
rect 40770 699864 40776 699916
rect 40828 699904 40834 699916
rect 465077 699907 465135 699913
rect 465077 699904 465089 699907
rect 40828 699876 465089 699904
rect 40828 699864 40834 699876
rect 465077 699873 465089 699876
rect 465123 699873 465135 699907
rect 465077 699867 465135 699873
rect 18690 699796 18696 699848
rect 18748 699836 18754 699848
rect 443825 699839 443883 699845
rect 443825 699836 443837 699839
rect 18748 699808 443837 699836
rect 18748 699796 18754 699808
rect 443825 699805 443837 699808
rect 443871 699805 443883 699839
rect 443825 699799 443883 699805
rect 14550 699728 14556 699780
rect 14608 699768 14614 699780
rect 440329 699771 440387 699777
rect 440329 699768 440341 699771
rect 14608 699740 440341 699768
rect 14608 699728 14614 699740
rect 440329 699737 440341 699740
rect 440375 699737 440387 699771
rect 440329 699731 440387 699737
rect 33870 699660 33876 699712
rect 33928 699700 33934 699712
rect 461489 699703 461547 699709
rect 461489 699700 461501 699703
rect 33928 699672 461501 699700
rect 33928 699660 33934 699672
rect 461489 699669 461501 699672
rect 461535 699669 461547 699703
rect 461489 699663 461547 699669
rect 349065 699635 349123 699641
rect 349065 699601 349077 699635
rect 349111 699632 349123 699635
rect 362129 699635 362187 699641
rect 362129 699632 362141 699635
rect 349111 699604 362141 699632
rect 349111 699601 349123 699604
rect 349065 699595 349123 699601
rect 362129 699601 362141 699604
rect 362175 699601 362187 699635
rect 362129 699595 362187 699601
rect 362221 699635 362279 699641
rect 362221 699601 362233 699635
rect 362267 699632 362279 699635
rect 369673 699635 369731 699641
rect 369673 699632 369685 699635
rect 362267 699604 369685 699632
rect 362267 699601 362279 699604
rect 362221 699595 362279 699601
rect 369673 699601 369685 699604
rect 369719 699601 369731 699635
rect 369673 699595 369731 699601
rect 369857 699635 369915 699641
rect 369857 699601 369869 699635
rect 369903 699632 369915 699635
rect 391109 699635 391167 699641
rect 391109 699632 391121 699635
rect 369903 699604 391121 699632
rect 369903 699601 369915 699604
rect 369857 699595 369915 699601
rect 391109 699601 391121 699604
rect 391155 699601 391167 699635
rect 401689 699635 401747 699641
rect 401689 699632 401701 699635
rect 391109 699595 391167 699601
rect 393286 699604 401701 699632
rect 363049 699567 363107 699573
rect 363049 699533 363061 699567
rect 363095 699564 363107 699567
rect 393286 699564 393314 699604
rect 401689 699601 401701 699604
rect 401735 699601 401747 699635
rect 401689 699595 401747 699601
rect 363095 699536 393314 699564
rect 363095 699533 363107 699536
rect 363049 699527 363107 699533
rect 3510 684428 3516 684480
rect 3568 684468 3574 684480
rect 182174 684468 182180 684480
rect 3568 684440 182180 684468
rect 3568 684428 3574 684440
rect 182174 684428 182180 684440
rect 182232 684428 182238 684480
rect 3050 671984 3056 672036
rect 3108 672024 3114 672036
rect 18690 672024 18696 672036
rect 3108 671996 18696 672024
rect 3108 671984 3114 671996
rect 18690 671984 18696 671996
rect 18748 671984 18754 672036
rect 3510 658180 3516 658232
rect 3568 658220 3574 658232
rect 14550 658220 14556 658232
rect 3568 658192 14556 658220
rect 3568 658180 3574 658192
rect 14550 658180 14556 658192
rect 14608 658180 14614 658232
rect 3234 633360 3240 633412
rect 3292 633400 3298 633412
rect 182266 633400 182272 633412
rect 3292 633372 182272 633400
rect 3292 633360 3298 633372
rect 182266 633360 182272 633372
rect 182324 633360 182330 633412
rect 3326 619556 3332 619608
rect 3384 619596 3390 619608
rect 35250 619596 35256 619608
rect 3384 619568 35256 619596
rect 3384 619556 3390 619568
rect 35250 619556 35256 619568
rect 35308 619556 35314 619608
rect 3234 607112 3240 607164
rect 3292 607152 3298 607164
rect 32490 607152 32496 607164
rect 3292 607124 32496 607152
rect 3292 607112 3298 607124
rect 32490 607112 32496 607124
rect 32548 607112 32554 607164
rect 3142 580932 3148 580984
rect 3200 580972 3206 580984
rect 182358 580972 182364 580984
rect 3200 580944 182364 580972
rect 3200 580932 3206 580944
rect 182358 580932 182364 580944
rect 182416 580932 182422 580984
rect 3510 567128 3516 567180
rect 3568 567168 3574 567180
rect 40770 567168 40776 567180
rect 3568 567140 40776 567168
rect 3568 567128 3574 567140
rect 40770 567128 40776 567140
rect 40828 567128 40834 567180
rect 3510 554684 3516 554736
rect 3568 554724 3574 554736
rect 33870 554724 33876 554736
rect 3568 554696 33876 554724
rect 3568 554684 3574 554696
rect 33870 554684 33876 554696
rect 33928 554684 33934 554736
rect 2866 528504 2872 528556
rect 2924 528544 2930 528556
rect 182450 528544 182456 528556
rect 2924 528516 182456 528544
rect 2924 528504 2930 528516
rect 182450 528504 182456 528516
rect 182508 528504 182514 528556
rect 3510 516060 3516 516112
rect 3568 516100 3574 516112
rect 18598 516100 18604 516112
rect 3568 516072 18604 516100
rect 3568 516060 3574 516072
rect 18598 516060 18604 516072
rect 18656 516060 18662 516112
rect 3510 502256 3516 502308
rect 3568 502296 3574 502308
rect 14458 502296 14464 502308
rect 3568 502268 14464 502296
rect 3568 502256 3574 502268
rect 14458 502256 14464 502268
rect 14516 502256 14522 502308
rect 3510 476008 3516 476060
rect 3568 476048 3574 476060
rect 182542 476048 182548 476060
rect 3568 476020 182548 476048
rect 3568 476008 3574 476020
rect 182542 476008 182548 476020
rect 182600 476008 182606 476060
rect 3234 463632 3240 463684
rect 3292 463672 3298 463684
rect 35158 463672 35164 463684
rect 3292 463644 35164 463672
rect 3292 463632 3298 463644
rect 35158 463632 35164 463644
rect 35216 463632 35222 463684
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 32398 449868 32404 449880
rect 3384 449840 32404 449868
rect 3384 449828 3390 449840
rect 32398 449828 32404 449840
rect 32456 449828 32462 449880
rect 3510 423580 3516 423632
rect 3568 423620 3574 423632
rect 182634 423620 182640 423632
rect 3568 423592 182640 423620
rect 3568 423580 3574 423592
rect 182634 423580 182640 423592
rect 182692 423580 182698 423632
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 25498 411244 25504 411256
rect 3016 411216 25504 411244
rect 3016 411204 3022 411216
rect 25498 411204 25504 411216
rect 25556 411204 25562 411256
rect 3234 398760 3240 398812
rect 3292 398800 3298 398812
rect 17218 398800 17224 398812
rect 3292 398772 17224 398800
rect 3292 398760 3298 398772
rect 17218 398760 17224 398772
rect 17276 398760 17282 398812
rect 3510 372512 3516 372564
rect 3568 372552 3574 372564
rect 182726 372552 182732 372564
rect 3568 372524 182732 372552
rect 3568 372512 3574 372524
rect 182726 372512 182732 372524
rect 182784 372512 182790 372564
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 29638 358748 29644 358760
rect 3384 358720 29644 358748
rect 3384 358708 3390 358720
rect 29638 358708 29644 358720
rect 29696 358708 29702 358760
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 177298 346372 177304 346384
rect 3200 346344 177304 346372
rect 3200 346332 3206 346344
rect 177298 346332 177304 346344
rect 177356 346332 177362 346384
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 182726 318832 182732 318844
rect 3384 318804 182732 318832
rect 3384 318792 3390 318804
rect 182726 318792 182732 318804
rect 182784 318792 182790 318844
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 33778 306320 33784 306332
rect 3568 306292 33784 306320
rect 3568 306280 3574 306292
rect 33778 306280 33784 306292
rect 33836 306280 33842 306332
rect 182818 302948 182824 303000
rect 182876 302988 182882 303000
rect 182876 302960 580304 302988
rect 182876 302948 182882 302960
rect 181806 302880 181812 302932
rect 181864 302920 181870 302932
rect 181864 302892 567194 302920
rect 181864 302880 181870 302892
rect 567166 302376 567194 302892
rect 580276 302456 580304 302960
rect 580258 302404 580264 302456
rect 580316 302404 580322 302456
rect 580350 302376 580356 302388
rect 567166 302348 580356 302376
rect 580350 302336 580356 302348
rect 580408 302336 580414 302388
rect 182174 299480 182180 299532
rect 182232 299520 182238 299532
rect 183186 299520 183192 299532
rect 182232 299492 183192 299520
rect 182232 299480 182238 299492
rect 183186 299480 183192 299492
rect 183244 299480 183250 299532
rect 183554 299480 183560 299532
rect 183612 299520 183618 299532
rect 184382 299520 184388 299532
rect 183612 299492 184388 299520
rect 183612 299480 183618 299492
rect 184382 299480 184388 299492
rect 184440 299480 184446 299532
rect 351914 299480 351920 299532
rect 351972 299520 351978 299532
rect 352374 299520 352380 299532
rect 351972 299492 352380 299520
rect 351972 299480 351978 299492
rect 352374 299480 352380 299492
rect 352432 299480 352438 299532
rect 353386 299480 353392 299532
rect 353444 299520 353450 299532
rect 354030 299520 354036 299532
rect 353444 299492 354036 299520
rect 353444 299480 353450 299492
rect 354030 299480 354036 299492
rect 354088 299480 354094 299532
rect 367094 299480 367100 299532
rect 367152 299520 367158 299532
rect 367830 299520 367836 299532
rect 367152 299492 367836 299520
rect 367152 299480 367158 299492
rect 367830 299480 367836 299492
rect 367888 299480 367894 299532
rect 440234 299480 440240 299532
rect 440292 299520 440298 299532
rect 440878 299520 440884 299532
rect 440292 299492 440884 299520
rect 440292 299480 440298 299492
rect 440878 299480 440884 299492
rect 440936 299480 440942 299532
rect 493229 299523 493287 299529
rect 493229 299489 493241 299523
rect 493275 299520 493287 299523
rect 493275 299492 494008 299520
rect 493275 299489 493287 299492
rect 493229 299483 493287 299489
rect 107562 299412 107568 299464
rect 107620 299452 107626 299464
rect 256142 299452 256148 299464
rect 107620 299424 256148 299452
rect 107620 299412 107626 299424
rect 256142 299412 256148 299424
rect 256200 299412 256206 299464
rect 258074 299412 258080 299464
rect 258132 299452 258138 299464
rect 265066 299452 265072 299464
rect 258132 299424 265072 299452
rect 258132 299412 258138 299424
rect 265066 299412 265072 299424
rect 265124 299412 265130 299464
rect 265161 299455 265219 299461
rect 265161 299421 265173 299455
rect 265207 299452 265219 299455
rect 293494 299452 293500 299464
rect 265207 299424 293500 299452
rect 265207 299421 265219 299424
rect 265161 299415 265219 299421
rect 293494 299412 293500 299424
rect 293552 299412 293558 299464
rect 296070 299412 296076 299464
rect 296128 299452 296134 299464
rect 312998 299452 313004 299464
rect 296128 299424 313004 299452
rect 296128 299412 296134 299424
rect 312998 299412 313004 299424
rect 313056 299412 313062 299464
rect 335354 299412 335360 299464
rect 335412 299452 335418 299464
rect 336182 299452 336188 299464
rect 335412 299424 336188 299452
rect 335412 299412 335418 299424
rect 336182 299412 336188 299424
rect 336240 299412 336246 299464
rect 338114 299412 338120 299464
rect 338172 299452 338178 299464
rect 338574 299452 338580 299464
rect 338172 299424 338580 299452
rect 338172 299412 338178 299424
rect 338574 299412 338580 299424
rect 338632 299412 338638 299464
rect 339494 299412 339500 299464
rect 339552 299452 339558 299464
rect 340230 299452 340236 299464
rect 339552 299424 340236 299452
rect 339552 299412 339558 299424
rect 340230 299412 340236 299424
rect 340288 299412 340294 299464
rect 340325 299455 340383 299461
rect 340325 299421 340337 299455
rect 340371 299452 340383 299455
rect 414382 299452 414388 299464
rect 340371 299424 414388 299452
rect 340371 299421 340383 299424
rect 340325 299415 340383 299421
rect 414382 299412 414388 299424
rect 414440 299412 414446 299464
rect 416682 299412 416688 299464
rect 416740 299452 416746 299464
rect 421561 299455 421619 299461
rect 416740 299424 421512 299452
rect 416740 299412 416746 299424
rect 103422 299344 103428 299396
rect 103480 299384 103486 299396
rect 253750 299384 253756 299396
rect 103480 299356 253756 299384
rect 103480 299344 103486 299356
rect 253750 299344 253756 299356
rect 253808 299344 253814 299396
rect 273162 299384 273168 299396
rect 253860 299356 273168 299384
rect 90358 299276 90364 299328
rect 90416 299316 90422 299328
rect 243998 299316 244004 299328
rect 90416 299288 244004 299316
rect 90416 299276 90422 299288
rect 243998 299276 244004 299288
rect 244056 299276 244062 299328
rect 246942 299276 246948 299328
rect 247000 299316 247006 299328
rect 248046 299316 248052 299328
rect 247000 299288 248052 299316
rect 247000 299276 247006 299288
rect 248046 299276 248052 299288
rect 248104 299276 248110 299328
rect 253290 299276 253296 299328
rect 253348 299316 253354 299328
rect 253860 299316 253888 299356
rect 273162 299344 273168 299356
rect 273220 299344 273226 299396
rect 274082 299344 274088 299396
rect 274140 299384 274146 299396
rect 317874 299384 317880 299396
rect 274140 299356 317880 299384
rect 274140 299344 274146 299356
rect 317874 299344 317880 299356
rect 317932 299344 317938 299396
rect 331858 299344 331864 299396
rect 331916 299384 331922 299396
rect 409506 299384 409512 299396
rect 331916 299356 409512 299384
rect 331916 299344 331922 299356
rect 409506 299344 409512 299356
rect 409564 299344 409570 299396
rect 410518 299344 410524 299396
rect 410576 299384 410582 299396
rect 416038 299384 416044 299396
rect 410576 299356 416044 299384
rect 410576 299344 410582 299356
rect 416038 299344 416044 299356
rect 416096 299344 416102 299396
rect 420914 299344 420920 299396
rect 420972 299384 420978 299396
rect 421374 299384 421380 299396
rect 420972 299356 421380 299384
rect 420972 299344 420978 299356
rect 421374 299344 421380 299356
rect 421432 299344 421438 299396
rect 421484 299384 421512 299424
rect 421561 299421 421573 299455
rect 421607 299452 421619 299455
rect 467098 299452 467104 299464
rect 421607 299424 467104 299452
rect 421607 299421 421619 299424
rect 421561 299415 421619 299421
rect 467098 299412 467104 299424
rect 467156 299412 467162 299464
rect 473998 299412 474004 299464
rect 474056 299452 474062 299464
rect 479334 299452 479340 299464
rect 474056 299424 479340 299452
rect 474056 299412 474062 299424
rect 479334 299412 479340 299424
rect 479392 299412 479398 299464
rect 479429 299455 479487 299461
rect 479429 299421 479441 299455
rect 479475 299452 479487 299455
rect 493870 299452 493876 299464
rect 479475 299424 493876 299452
rect 479475 299421 479487 299424
rect 479429 299415 479487 299421
rect 493870 299412 493876 299424
rect 493928 299412 493934 299464
rect 493980 299452 494008 299492
rect 501230 299452 501236 299464
rect 493980 299424 501236 299452
rect 501230 299412 501236 299424
rect 501288 299412 501294 299464
rect 501509 299455 501567 299461
rect 501509 299421 501521 299455
rect 501555 299452 501567 299455
rect 523126 299452 523132 299464
rect 501555 299424 523132 299452
rect 501555 299421 501567 299424
rect 501509 299415 501567 299421
rect 523126 299412 523132 299424
rect 523184 299412 523190 299464
rect 526438 299412 526444 299464
rect 526496 299452 526502 299464
rect 541802 299452 541808 299464
rect 526496 299424 541808 299452
rect 526496 299412 526502 299424
rect 541802 299412 541808 299424
rect 541860 299412 541866 299464
rect 547138 299412 547144 299464
rect 547196 299452 547202 299464
rect 557166 299452 557172 299464
rect 547196 299424 557172 299452
rect 547196 299412 547202 299424
rect 557166 299412 557172 299424
rect 557224 299412 557230 299464
rect 467926 299384 467932 299396
rect 421484 299356 467932 299384
rect 467926 299344 467932 299356
rect 467984 299344 467990 299396
rect 468036 299356 470594 299384
rect 253348 299288 253888 299316
rect 253937 299319 253995 299325
rect 253348 299276 253354 299288
rect 253937 299285 253949 299319
rect 253983 299316 253995 299319
rect 298370 299316 298376 299328
rect 253983 299288 298376 299316
rect 253983 299285 253995 299288
rect 253937 299279 253995 299285
rect 298370 299276 298376 299288
rect 298428 299276 298434 299328
rect 300118 299276 300124 299328
rect 300176 299316 300182 299328
rect 300857 299319 300915 299325
rect 300857 299316 300869 299319
rect 300176 299288 300869 299316
rect 300176 299276 300182 299288
rect 300857 299285 300869 299288
rect 300903 299285 300915 299319
rect 300857 299279 300915 299285
rect 300949 299319 301007 299325
rect 300949 299285 300961 299319
rect 300995 299316 301007 299319
rect 308122 299316 308128 299328
rect 300995 299288 308128 299316
rect 300995 299285 301007 299288
rect 300949 299279 301007 299285
rect 308122 299276 308128 299288
rect 308180 299276 308186 299328
rect 313274 299276 313280 299328
rect 313332 299316 313338 299328
rect 314286 299316 314292 299328
rect 313332 299288 314292 299316
rect 313332 299276 313338 299288
rect 314286 299276 314292 299288
rect 314344 299276 314350 299328
rect 320174 299276 320180 299328
rect 320232 299316 320238 299328
rect 320726 299316 320732 299328
rect 320232 299288 320732 299316
rect 320232 299276 320238 299288
rect 320726 299276 320732 299288
rect 320784 299276 320790 299328
rect 325694 299276 325700 299328
rect 325752 299316 325758 299328
rect 326430 299316 326436 299328
rect 325752 299288 326436 299316
rect 325752 299276 325758 299288
rect 326430 299276 326436 299288
rect 326488 299276 326494 299328
rect 327718 299276 327724 299328
rect 327776 299316 327782 299328
rect 404630 299316 404636 299328
rect 327776 299288 404636 299316
rect 327776 299276 327782 299288
rect 404630 299276 404636 299288
rect 404688 299276 404694 299328
rect 408402 299276 408408 299328
rect 408460 299316 408466 299328
rect 463050 299316 463056 299328
rect 408460 299288 463056 299316
rect 408460 299276 408466 299288
rect 463050 299276 463056 299288
rect 463108 299276 463114 299328
rect 467742 299276 467748 299328
rect 467800 299316 467806 299328
rect 468036 299316 468064 299356
rect 467800 299288 468064 299316
rect 467800 299276 467806 299288
rect 469214 299276 469220 299328
rect 469272 299316 469278 299328
rect 470134 299316 470140 299328
rect 469272 299288 470140 299316
rect 469272 299276 469278 299288
rect 470134 299276 470140 299288
rect 470192 299276 470198 299328
rect 470566 299316 470594 299356
rect 472618 299344 472624 299396
rect 472676 299384 472682 299396
rect 476850 299384 476856 299396
rect 472676 299356 476856 299384
rect 472676 299344 472682 299356
rect 476850 299344 476856 299356
rect 476908 299344 476914 299396
rect 478138 299344 478144 299396
rect 478196 299384 478202 299396
rect 506106 299384 506112 299396
rect 478196 299356 506112 299384
rect 478196 299344 478202 299356
rect 506106 299344 506112 299356
rect 506164 299344 506170 299396
rect 507762 299344 507768 299396
rect 507820 299384 507826 299396
rect 530394 299384 530400 299396
rect 507820 299356 530400 299384
rect 507820 299344 507826 299356
rect 530394 299344 530400 299356
rect 530452 299344 530458 299396
rect 530578 299344 530584 299396
rect 530636 299384 530642 299396
rect 536098 299384 536104 299396
rect 530636 299356 536104 299384
rect 530636 299344 530642 299356
rect 536098 299344 536104 299356
rect 536156 299344 536162 299396
rect 549070 299384 549076 299396
rect 536208 299356 549076 299384
rect 503622 299316 503628 299328
rect 470566 299288 503628 299316
rect 503622 299276 503628 299288
rect 503680 299276 503686 299328
rect 504358 299276 504364 299328
rect 504416 299316 504422 299328
rect 506842 299316 506848 299328
rect 504416 299288 506848 299316
rect 504416 299276 504422 299288
rect 506842 299276 506848 299288
rect 506900 299276 506906 299328
rect 506937 299319 506995 299325
rect 506937 299285 506949 299319
rect 506983 299316 506995 299319
rect 522301 299319 522359 299325
rect 522301 299316 522313 299319
rect 506983 299288 522313 299316
rect 506983 299285 506995 299288
rect 506937 299279 506995 299285
rect 522301 299285 522313 299288
rect 522347 299285 522359 299319
rect 522301 299279 522359 299285
rect 522390 299276 522396 299328
rect 522448 299316 522454 299328
rect 524690 299316 524696 299328
rect 522448 299288 524696 299316
rect 522448 299276 522454 299288
rect 524690 299276 524696 299288
rect 524748 299276 524754 299328
rect 525150 299276 525156 299328
rect 525208 299316 525214 299328
rect 527174 299316 527180 299328
rect 525208 299288 527180 299316
rect 525208 299276 525214 299288
rect 527174 299276 527180 299288
rect 527232 299276 527238 299328
rect 529290 299276 529296 299328
rect 529348 299316 529354 299328
rect 531222 299316 531228 299328
rect 529348 299288 531228 299316
rect 529348 299276 529354 299288
rect 531222 299276 531228 299288
rect 531280 299276 531286 299328
rect 533982 299276 533988 299328
rect 534040 299316 534046 299328
rect 536208 299316 536236 299356
rect 549070 299344 549076 299356
rect 549128 299344 549134 299396
rect 558178 299344 558184 299396
rect 558236 299384 558242 299396
rect 565262 299384 565268 299396
rect 558236 299356 565268 299384
rect 558236 299344 558242 299356
rect 565262 299344 565268 299356
rect 565320 299344 565326 299396
rect 569218 299344 569224 299396
rect 569276 299384 569282 299396
rect 572622 299384 572628 299396
rect 569276 299356 572628 299384
rect 569276 299344 569282 299356
rect 572622 299344 572628 299356
rect 572680 299344 572686 299396
rect 534040 299288 536236 299316
rect 536285 299319 536343 299325
rect 534040 299276 534046 299288
rect 536285 299285 536297 299319
rect 536331 299316 536343 299319
rect 546678 299316 546684 299328
rect 536331 299288 546684 299316
rect 536331 299285 536343 299288
rect 536285 299279 536343 299285
rect 546678 299276 546684 299288
rect 546736 299276 546742 299328
rect 548518 299276 548524 299328
rect 548576 299316 548582 299328
rect 557994 299316 558000 299328
rect 548576 299288 558000 299316
rect 548576 299276 548582 299288
rect 557994 299276 558000 299288
rect 558052 299276 558058 299328
rect 560938 299276 560944 299328
rect 560996 299316 561002 299328
rect 566918 299316 566924 299328
rect 560996 299288 566924 299316
rect 560996 299276 561002 299288
rect 566918 299276 566924 299288
rect 566976 299276 566982 299328
rect 574002 299276 574008 299328
rect 574060 299316 574066 299328
rect 575842 299316 575848 299328
rect 574060 299288 575848 299316
rect 574060 299276 574066 299288
rect 575842 299276 575848 299288
rect 575900 299276 575906 299328
rect 582374 299276 582380 299328
rect 582432 299316 582438 299328
rect 583113 299319 583171 299325
rect 583113 299316 583125 299319
rect 582432 299288 583125 299316
rect 582432 299276 582438 299288
rect 583113 299285 583125 299288
rect 583159 299285 583171 299319
rect 583113 299279 583171 299285
rect 50338 299208 50344 299260
rect 50396 299248 50402 299260
rect 214742 299248 214748 299260
rect 50396 299220 214748 299248
rect 50396 299208 50402 299220
rect 214742 299208 214748 299220
rect 214800 299208 214806 299260
rect 232498 299208 232504 299260
rect 232556 299248 232562 299260
rect 263502 299248 263508 299260
rect 232556 299220 263508 299248
rect 232556 299208 232562 299220
rect 263502 299208 263508 299220
rect 263560 299208 263566 299260
rect 263686 299208 263692 299260
rect 263744 299248 263750 299260
rect 274818 299248 274824 299260
rect 263744 299220 274824 299248
rect 263744 299208 263750 299220
rect 274818 299208 274824 299220
rect 274876 299208 274882 299260
rect 281350 299208 281356 299260
rect 281408 299248 281414 299260
rect 283742 299248 283748 299260
rect 281408 299220 283748 299248
rect 281408 299208 281414 299220
rect 283742 299208 283748 299220
rect 283800 299208 283806 299260
rect 285674 299208 285680 299260
rect 285732 299248 285738 299260
rect 286686 299248 286692 299260
rect 285732 299220 286692 299248
rect 285732 299208 285738 299220
rect 286686 299208 286692 299220
rect 286744 299208 286750 299260
rect 286781 299251 286839 299257
rect 286781 299217 286793 299251
rect 286827 299248 286839 299251
rect 355962 299248 355968 299260
rect 286827 299220 355968 299248
rect 286827 299217 286839 299220
rect 286781 299211 286839 299217
rect 355962 299208 355968 299220
rect 356020 299208 356026 299260
rect 357434 299208 357440 299260
rect 357492 299248 357498 299260
rect 358078 299248 358084 299260
rect 357492 299220 358084 299248
rect 357492 299208 357498 299220
rect 358078 299208 358084 299220
rect 358136 299208 358142 299260
rect 358814 299208 358820 299260
rect 358872 299248 358878 299260
rect 359734 299248 359740 299260
rect 358872 299220 359740 299248
rect 358872 299208 358878 299220
rect 359734 299208 359740 299220
rect 359792 299208 359798 299260
rect 362218 299208 362224 299260
rect 362276 299248 362282 299260
rect 363230 299248 363236 299260
rect 362276 299220 363236 299248
rect 362276 299208 362282 299220
rect 363230 299208 363236 299220
rect 363288 299208 363294 299260
rect 363325 299251 363383 299257
rect 363325 299217 363337 299251
rect 363371 299248 363383 299251
rect 429010 299248 429016 299260
rect 363371 299220 429016 299248
rect 363371 299217 363383 299220
rect 363325 299211 363383 299217
rect 429010 299208 429016 299220
rect 429068 299208 429074 299260
rect 430574 299208 430580 299260
rect 430632 299248 430638 299260
rect 431126 299248 431132 299260
rect 430632 299220 431132 299248
rect 430632 299208 430638 299220
rect 431126 299208 431132 299220
rect 431184 299208 431190 299260
rect 431221 299251 431279 299257
rect 431221 299217 431233 299251
rect 431267 299248 431279 299251
rect 477678 299248 477684 299260
rect 431267 299220 477684 299248
rect 431267 299217 431279 299220
rect 431221 299211 431279 299217
rect 477678 299208 477684 299220
rect 477736 299208 477742 299260
rect 478230 299208 478236 299260
rect 478288 299248 478294 299260
rect 480070 299248 480076 299260
rect 478288 299220 480076 299248
rect 478288 299208 478294 299220
rect 480070 299208 480076 299220
rect 480128 299208 480134 299260
rect 480162 299208 480168 299260
rect 480220 299248 480226 299260
rect 484946 299248 484952 299260
rect 480220 299220 484952 299248
rect 480220 299208 480226 299220
rect 484946 299208 484952 299220
rect 485004 299208 485010 299260
rect 491113 299251 491171 299257
rect 491113 299217 491125 299251
rect 491159 299248 491171 299251
rect 493229 299251 493287 299257
rect 493229 299248 493241 299251
rect 491159 299220 493241 299248
rect 491159 299217 491171 299220
rect 491113 299211 491171 299217
rect 493229 299217 493241 299220
rect 493275 299217 493287 299251
rect 493229 299211 493287 299217
rect 493318 299208 493324 299260
rect 493376 299248 493382 299260
rect 496354 299248 496360 299260
rect 493376 299220 496360 299248
rect 493376 299208 493382 299220
rect 496354 299208 496360 299220
rect 496412 299208 496418 299260
rect 496449 299251 496507 299257
rect 496449 299217 496461 299251
rect 496495 299248 496507 299251
rect 519078 299248 519084 299260
rect 496495 299220 519084 299248
rect 496495 299217 496507 299220
rect 496449 299211 496507 299217
rect 519078 299208 519084 299220
rect 519136 299208 519142 299260
rect 519538 299208 519544 299260
rect 519596 299248 519602 299260
rect 523954 299248 523960 299260
rect 519596 299220 523960 299248
rect 519596 299208 519602 299220
rect 523954 299208 523960 299220
rect 524012 299208 524018 299260
rect 524049 299251 524107 299257
rect 524049 299217 524061 299251
rect 524095 299248 524107 299251
rect 539318 299248 539324 299260
rect 524095 299220 539324 299248
rect 524095 299217 524107 299220
rect 524049 299211 524107 299217
rect 539318 299208 539324 299220
rect 539376 299208 539382 299260
rect 540238 299208 540244 299260
rect 540296 299248 540302 299260
rect 550726 299248 550732 299260
rect 540296 299220 550732 299248
rect 540296 299208 540302 299220
rect 550726 299208 550732 299220
rect 550784 299208 550790 299260
rect 551922 299208 551928 299260
rect 551980 299248 551986 299260
rect 561214 299248 561220 299260
rect 551980 299220 561220 299248
rect 551980 299208 551986 299220
rect 561214 299208 561220 299220
rect 561272 299208 561278 299260
rect 572622 299208 572628 299260
rect 572680 299248 572686 299260
rect 575014 299248 575020 299260
rect 572680 299220 575020 299248
rect 572680 299208 572686 299220
rect 575014 299208 575020 299220
rect 575072 299208 575078 299260
rect 35158 299140 35164 299192
rect 35216 299180 35222 299192
rect 194873 299183 194931 299189
rect 194873 299180 194885 299183
rect 35216 299152 194885 299180
rect 35216 299140 35222 299152
rect 194873 299149 194885 299152
rect 194919 299149 194931 299183
rect 194873 299143 194931 299149
rect 195974 299140 195980 299192
rect 196032 299180 196038 299192
rect 196526 299180 196532 299192
rect 196032 299152 196532 299180
rect 196032 299140 196038 299152
rect 196526 299140 196532 299152
rect 196584 299140 196590 299192
rect 201494 299140 201500 299192
rect 201552 299180 201558 299192
rect 202230 299180 202236 299192
rect 201552 299152 202236 299180
rect 201552 299140 201558 299152
rect 202230 299140 202236 299152
rect 202288 299140 202294 299192
rect 220078 299140 220084 299192
rect 220136 299180 220142 299192
rect 241606 299180 241612 299192
rect 220136 299152 241612 299180
rect 220136 299140 220142 299152
rect 241606 299140 241612 299152
rect 241664 299140 241670 299192
rect 246482 299140 246488 299192
rect 246540 299180 246546 299192
rect 300762 299180 300768 299192
rect 246540 299152 300768 299180
rect 246540 299140 246546 299152
rect 300762 299140 300768 299152
rect 300820 299140 300826 299192
rect 300857 299183 300915 299189
rect 300857 299149 300869 299183
rect 300903 299180 300915 299183
rect 312170 299180 312176 299192
rect 300903 299152 312176 299180
rect 300903 299149 300915 299152
rect 300857 299143 300915 299149
rect 312170 299140 312176 299152
rect 312228 299140 312234 299192
rect 312538 299140 312544 299192
rect 312596 299180 312602 299192
rect 319438 299180 319444 299192
rect 312596 299152 319444 299180
rect 312596 299140 312602 299152
rect 319438 299140 319444 299152
rect 319496 299140 319502 299192
rect 322198 299140 322204 299192
rect 322256 299180 322262 299192
rect 399386 299180 399392 299192
rect 322256 299152 399392 299180
rect 322256 299140 322262 299152
rect 399386 299140 399392 299152
rect 399444 299140 399450 299192
rect 399478 299140 399484 299192
rect 399536 299180 399542 299192
rect 402238 299180 402244 299192
rect 399536 299152 402244 299180
rect 399536 299140 399542 299152
rect 402238 299140 402244 299152
rect 402296 299140 402302 299192
rect 402333 299183 402391 299189
rect 402333 299149 402345 299183
rect 402379 299180 402391 299183
rect 454313 299183 454371 299189
rect 454313 299180 454325 299183
rect 402379 299152 454325 299180
rect 402379 299149 402391 299152
rect 402333 299143 402391 299149
rect 454313 299149 454325 299152
rect 454359 299149 454371 299183
rect 454313 299143 454371 299149
rect 456058 299140 456064 299192
rect 456116 299180 456122 299192
rect 460658 299180 460664 299192
rect 456116 299152 460664 299180
rect 456116 299140 456122 299152
rect 460658 299140 460664 299152
rect 460716 299140 460722 299192
rect 460753 299183 460811 299189
rect 460753 299149 460765 299183
rect 460799 299180 460811 299183
rect 497182 299180 497188 299192
rect 460799 299152 497188 299180
rect 460799 299149 460811 299152
rect 460753 299143 460811 299149
rect 497182 299140 497188 299152
rect 497240 299140 497246 299192
rect 503622 299140 503628 299192
rect 503680 299180 503686 299192
rect 506937 299183 506995 299189
rect 506937 299180 506949 299183
rect 503680 299152 506949 299180
rect 503680 299140 503686 299152
rect 506937 299149 506949 299152
rect 506983 299149 506995 299183
rect 506937 299143 506995 299149
rect 507029 299183 507087 299189
rect 507029 299149 507041 299183
rect 507075 299180 507087 299183
rect 526346 299180 526352 299192
rect 507075 299152 526352 299180
rect 507075 299149 507087 299152
rect 507029 299143 507087 299149
rect 526346 299140 526352 299152
rect 526404 299140 526410 299192
rect 527082 299140 527088 299192
rect 527140 299180 527146 299192
rect 544194 299180 544200 299192
rect 527140 299152 544200 299180
rect 527140 299140 527146 299152
rect 544194 299140 544200 299152
rect 544252 299140 544258 299192
rect 544378 299140 544384 299192
rect 544436 299180 544442 299192
rect 555326 299180 555332 299192
rect 544436 299152 555332 299180
rect 544436 299140 544442 299152
rect 555326 299140 555332 299152
rect 555384 299140 555390 299192
rect 555418 299140 555424 299192
rect 555476 299180 555482 299192
rect 562042 299180 562048 299192
rect 555476 299152 562048 299180
rect 555476 299140 555482 299152
rect 562042 299140 562048 299152
rect 562100 299140 562106 299192
rect 43438 299072 43444 299124
rect 43496 299112 43502 299124
rect 209958 299112 209964 299124
rect 43496 299084 209964 299112
rect 43496 299072 43502 299084
rect 209958 299072 209964 299084
rect 210016 299072 210022 299124
rect 217318 299072 217324 299124
rect 217376 299112 217382 299124
rect 239122 299112 239128 299124
rect 217376 299084 239128 299112
rect 217376 299072 217382 299084
rect 239122 299072 239128 299084
rect 239180 299072 239186 299124
rect 253198 299072 253204 299124
rect 253256 299112 253262 299124
rect 295886 299112 295892 299124
rect 253256 299084 295892 299112
rect 253256 299072 253262 299084
rect 295886 299072 295892 299084
rect 295944 299072 295950 299124
rect 295978 299072 295984 299124
rect 296036 299112 296042 299124
rect 296036 299084 376708 299112
rect 296036 299072 296042 299084
rect 33778 299004 33784 299056
rect 33836 299044 33842 299056
rect 205082 299044 205088 299056
rect 33836 299016 205088 299044
rect 33836 299004 33842 299016
rect 205082 299004 205088 299016
rect 205140 299004 205146 299056
rect 227070 299004 227076 299056
rect 227128 299044 227134 299056
rect 258626 299044 258632 299056
rect 227128 299016 258632 299044
rect 227128 299004 227134 299016
rect 258626 299004 258632 299016
rect 258684 299004 258690 299056
rect 262858 299004 262864 299056
rect 262916 299044 262922 299056
rect 279694 299044 279700 299056
rect 262916 299016 279700 299044
rect 262916 299004 262922 299016
rect 279694 299004 279700 299016
rect 279752 299004 279758 299056
rect 282178 299004 282184 299056
rect 282236 299044 282242 299056
rect 370590 299044 370596 299056
rect 282236 299016 370596 299044
rect 282236 299004 282242 299016
rect 370590 299004 370596 299016
rect 370648 299004 370654 299056
rect 371878 299004 371884 299056
rect 371936 299044 371942 299056
rect 372982 299044 372988 299056
rect 371936 299016 372988 299044
rect 371936 299004 371942 299016
rect 372982 299004 372988 299016
rect 373040 299004 373046 299056
rect 373902 299004 373908 299056
rect 373960 299044 373966 299056
rect 376481 299047 376539 299053
rect 376481 299044 376493 299047
rect 373960 299016 376493 299044
rect 373960 299004 373966 299016
rect 376481 299013 376493 299016
rect 376527 299013 376539 299047
rect 376481 299007 376539 299013
rect 29638 298936 29644 298988
rect 29696 298976 29702 298988
rect 200206 298976 200212 298988
rect 29696 298948 200212 298976
rect 29696 298936 29702 298948
rect 200206 298936 200212 298948
rect 200264 298936 200270 298988
rect 214558 298936 214564 298988
rect 214616 298976 214622 298988
rect 234246 298976 234252 298988
rect 214616 298948 234252 298976
rect 214616 298936 214622 298948
rect 234246 298936 234252 298948
rect 234304 298936 234310 298988
rect 234522 298936 234528 298988
rect 234580 298976 234586 298988
rect 268378 298976 268384 298988
rect 234580 298948 268384 298976
rect 234580 298936 234586 298948
rect 268378 298936 268384 298948
rect 268436 298936 268442 298988
rect 268838 298936 268844 298988
rect 268896 298976 268902 298988
rect 280982 298976 280988 298988
rect 268896 298948 280988 298976
rect 268896 298936 268902 298948
rect 280982 298936 280988 298948
rect 281040 298936 281046 298988
rect 284938 298936 284944 298988
rect 284996 298976 285002 298988
rect 375466 298976 375472 298988
rect 284996 298948 375472 298976
rect 284996 298936 285002 298948
rect 375466 298936 375472 298948
rect 375524 298936 375530 298988
rect 376680 298976 376708 299084
rect 376754 299072 376760 299124
rect 376812 299112 376818 299124
rect 377582 299112 377588 299124
rect 376812 299084 377588 299112
rect 376812 299072 376818 299084
rect 377582 299072 377588 299084
rect 377640 299072 377646 299124
rect 380158 299072 380164 299124
rect 380216 299112 380222 299124
rect 442810 299112 442816 299124
rect 380216 299084 442816 299112
rect 380216 299072 380222 299084
rect 442810 299072 442816 299084
rect 442868 299072 442874 299124
rect 443638 299072 443644 299124
rect 443696 299112 443702 299124
rect 445202 299112 445208 299124
rect 443696 299084 445208 299112
rect 443696 299072 443702 299084
rect 445202 299072 445208 299084
rect 445260 299072 445266 299124
rect 449158 299072 449164 299124
rect 449216 299112 449222 299124
rect 450078 299112 450084 299124
rect 449216 299084 450084 299112
rect 449216 299072 449222 299084
rect 450078 299072 450084 299084
rect 450136 299072 450142 299124
rect 450173 299115 450231 299121
rect 450173 299081 450185 299115
rect 450219 299112 450231 299115
rect 491478 299112 491484 299124
rect 450219 299084 491484 299112
rect 450219 299081 450231 299084
rect 450173 299075 450231 299081
rect 491478 299072 491484 299084
rect 491536 299072 491542 299124
rect 493962 299072 493968 299124
rect 494020 299112 494026 299124
rect 521470 299112 521476 299124
rect 494020 299084 521476 299112
rect 494020 299072 494026 299084
rect 521470 299072 521476 299084
rect 521528 299072 521534 299124
rect 522301 299115 522359 299121
rect 522301 299081 522313 299115
rect 522347 299112 522359 299115
rect 528002 299112 528008 299124
rect 522347 299084 528008 299112
rect 522347 299081 522359 299084
rect 522301 299075 522359 299081
rect 528002 299072 528008 299084
rect 528060 299072 528066 299124
rect 528097 299115 528155 299121
rect 528097 299081 528109 299115
rect 528143 299112 528155 299115
rect 540146 299112 540152 299124
rect 528143 299084 540152 299112
rect 528143 299081 528155 299084
rect 528097 299075 528155 299081
rect 540146 299072 540152 299084
rect 540204 299072 540210 299124
rect 543366 299112 543372 299124
rect 540808 299084 543372 299112
rect 376849 299047 376907 299053
rect 376849 299013 376861 299047
rect 376895 299044 376907 299047
rect 435269 299047 435327 299053
rect 435269 299044 435281 299047
rect 376895 299016 435281 299044
rect 376895 299013 376907 299016
rect 376849 299007 376907 299013
rect 435269 299013 435281 299016
rect 435315 299013 435327 299047
rect 435269 299007 435327 299013
rect 435358 299004 435364 299056
rect 435416 299044 435422 299056
rect 436278 299044 436284 299056
rect 435416 299016 436284 299044
rect 435416 299004 435422 299016
rect 436278 299004 436284 299016
rect 436336 299004 436342 299056
rect 436738 299004 436744 299056
rect 436796 299044 436802 299056
rect 437934 299044 437940 299056
rect 436796 299016 437940 299044
rect 436796 299004 436802 299016
rect 437934 299004 437940 299016
rect 437992 299004 437998 299056
rect 438118 299004 438124 299056
rect 438176 299044 438182 299056
rect 482554 299044 482560 299056
rect 438176 299016 482560 299044
rect 438176 299004 438182 299016
rect 482554 299004 482560 299016
rect 482612 299004 482618 299056
rect 485682 299004 485688 299056
rect 485740 299044 485746 299056
rect 515306 299044 515312 299056
rect 485740 299016 515312 299044
rect 485740 299004 485746 299016
rect 515306 299004 515312 299016
rect 515364 299004 515370 299056
rect 515398 299004 515404 299056
rect 515456 299044 515462 299056
rect 535270 299044 535276 299056
rect 515456 299016 535276 299044
rect 515456 299004 515462 299016
rect 535270 299004 535276 299016
rect 535328 299004 535334 299056
rect 536190 299004 536196 299056
rect 536248 299044 536254 299056
rect 540808 299044 540836 299084
rect 543366 299072 543372 299084
rect 543424 299072 543430 299124
rect 545022 299072 545028 299124
rect 545080 299112 545086 299124
rect 556338 299112 556344 299124
rect 545080 299084 556344 299112
rect 545080 299072 545086 299084
rect 556338 299072 556344 299084
rect 556396 299072 556402 299124
rect 536248 299016 540836 299044
rect 536248 299004 536254 299016
rect 542998 299004 543004 299056
rect 543056 299044 543062 299056
rect 554774 299044 554780 299056
rect 543056 299016 554780 299044
rect 543056 299004 543062 299016
rect 554774 299004 554780 299016
rect 554832 299004 554838 299056
rect 380342 298976 380348 298988
rect 376680 298948 380348 298976
rect 380342 298936 380348 298948
rect 380400 298936 380406 298988
rect 380802 298936 380808 298988
rect 380860 298976 380866 298988
rect 442169 298979 442227 298985
rect 442169 298976 442181 298979
rect 380860 298948 442181 298976
rect 380860 298936 380866 298948
rect 442169 298945 442181 298948
rect 442215 298945 442227 298979
rect 442169 298939 442227 298945
rect 442258 298936 442264 298988
rect 442316 298976 442322 298988
rect 446030 298976 446036 298988
rect 442316 298948 446036 298976
rect 442316 298936 442322 298948
rect 446030 298936 446036 298948
rect 446088 298936 446094 298988
rect 449802 298936 449808 298988
rect 449860 298976 449866 298988
rect 450173 298979 450231 298985
rect 450173 298976 450185 298979
rect 449860 298948 450185 298976
rect 449860 298936 449866 298948
rect 450173 298945 450185 298948
rect 450219 298945 450231 298979
rect 450173 298939 450231 298945
rect 450265 298979 450323 298985
rect 450265 298945 450277 298979
rect 450311 298976 450323 298979
rect 487430 298976 487436 298988
rect 450311 298948 487436 298976
rect 450311 298945 450323 298948
rect 450265 298939 450323 298945
rect 487430 298936 487436 298948
rect 487488 298936 487494 298988
rect 489822 298936 489828 298988
rect 489880 298976 489886 298988
rect 518250 298976 518256 298988
rect 489880 298948 518256 298976
rect 489880 298936 489886 298948
rect 518250 298936 518256 298948
rect 518308 298936 518314 298988
rect 518802 298936 518808 298988
rect 518860 298976 518866 298988
rect 538490 298976 538496 298988
rect 518860 298948 538496 298976
rect 518860 298936 518866 298948
rect 538490 298936 538496 298948
rect 538548 298936 538554 298988
rect 540882 298936 540888 298988
rect 540940 298976 540946 298988
rect 553946 298976 553952 298988
rect 540940 298948 553952 298976
rect 540940 298936 540946 298948
rect 553946 298936 553952 298948
rect 554004 298936 554010 298988
rect 556798 298936 556804 298988
rect 556856 298976 556862 298988
rect 563698 298976 563704 298988
rect 556856 298948 563704 298976
rect 556856 298936 556862 298948
rect 563698 298936 563704 298948
rect 563756 298936 563762 298988
rect 18598 298868 18604 298920
rect 18656 298908 18662 298920
rect 192846 298908 192852 298920
rect 18656 298880 192852 298908
rect 18656 298868 18662 298880
rect 192846 298868 192852 298880
rect 192904 298868 192910 298920
rect 194873 298911 194931 298917
rect 194873 298877 194885 298911
rect 194919 298908 194931 298911
rect 199378 298908 199384 298920
rect 194919 298880 199384 298908
rect 194919 298877 194931 298880
rect 194873 298871 194931 298877
rect 199378 298868 199384 298880
rect 199436 298868 199442 298920
rect 211798 298868 211804 298920
rect 211856 298908 211862 298920
rect 224494 298908 224500 298920
rect 211856 298880 224500 298908
rect 211856 298868 211862 298880
rect 224494 298868 224500 298880
rect 224552 298868 224558 298920
rect 251266 298908 251272 298920
rect 224604 298880 251272 298908
rect 17218 298800 17224 298852
rect 17276 298840 17282 298852
rect 193674 298840 193680 298852
rect 17276 298812 193680 298840
rect 17276 298800 17282 298812
rect 193674 298800 193680 298812
rect 193732 298800 193738 298852
rect 210418 298800 210424 298852
rect 210476 298840 210482 298852
rect 219618 298840 219624 298852
rect 210476 298812 219624 298840
rect 210476 298800 210482 298812
rect 219618 298800 219624 298812
rect 219676 298800 219682 298852
rect 224218 298800 224224 298852
rect 224276 298840 224282 298852
rect 224604 298840 224632 298880
rect 251266 298868 251272 298880
rect 251324 298868 251330 298920
rect 255958 298868 255964 298920
rect 256016 298908 256022 298920
rect 256016 298880 346992 298908
rect 256016 298868 256022 298880
rect 224276 298812 224632 298840
rect 224681 298843 224739 298849
rect 224276 298800 224282 298812
rect 224681 298809 224693 298843
rect 224727 298840 224739 298843
rect 246390 298840 246396 298852
rect 224727 298812 246396 298840
rect 224727 298809 224739 298812
rect 224681 298803 224739 298809
rect 246390 298800 246396 298812
rect 246448 298800 246454 298852
rect 249058 298800 249064 298852
rect 249116 298840 249122 298852
rect 346210 298840 346216 298852
rect 249116 298812 346216 298840
rect 249116 298800 249122 298812
rect 346210 298800 346216 298812
rect 346268 298800 346274 298852
rect 346964 298840 346992 298880
rect 347038 298868 347044 298920
rect 347096 298908 347102 298920
rect 348694 298908 348700 298920
rect 347096 298880 348700 298908
rect 347096 298868 347102 298880
rect 348694 298868 348700 298880
rect 348752 298868 348758 298920
rect 351822 298868 351828 298920
rect 351880 298908 351886 298920
rect 424134 298908 424140 298920
rect 351880 298880 424140 298908
rect 351880 298868 351886 298880
rect 424134 298868 424140 298880
rect 424192 298868 424198 298920
rect 430482 298868 430488 298920
rect 430540 298908 430546 298920
rect 431221 298911 431279 298917
rect 431221 298908 431233 298911
rect 430540 298880 431233 298908
rect 430540 298868 430546 298880
rect 431221 298877 431233 298880
rect 431267 298877 431279 298911
rect 474458 298908 474464 298920
rect 431221 298871 431279 298877
rect 431328 298880 474464 298908
rect 351086 298840 351092 298852
rect 346964 298812 351092 298840
rect 351086 298800 351092 298812
rect 351144 298800 351150 298852
rect 351181 298843 351239 298849
rect 351181 298809 351193 298843
rect 351227 298840 351239 298843
rect 419258 298840 419264 298852
rect 351227 298812 419264 298840
rect 351227 298809 351239 298812
rect 351181 298803 351239 298809
rect 419258 298800 419264 298812
rect 419316 298800 419322 298852
rect 424962 298800 424968 298852
rect 425020 298840 425026 298852
rect 431328 298840 431356 298880
rect 474458 298868 474464 298880
rect 474516 298868 474522 298920
rect 476758 298868 476764 298920
rect 476816 298908 476822 298920
rect 486602 298908 486608 298920
rect 476816 298880 486608 298908
rect 476816 298868 476822 298880
rect 486602 298868 486608 298880
rect 486660 298868 486666 298920
rect 487062 298868 487068 298920
rect 487120 298908 487126 298920
rect 516594 298908 516600 298920
rect 487120 298880 516600 298908
rect 487120 298868 487126 298880
rect 516594 298868 516600 298880
rect 516652 298868 516658 298920
rect 517422 298868 517428 298920
rect 517480 298908 517486 298920
rect 531133 298911 531191 298917
rect 531133 298908 531145 298911
rect 517480 298880 531145 298908
rect 517480 298868 517486 298880
rect 531133 298877 531145 298880
rect 531179 298877 531191 298911
rect 531133 298871 531191 298877
rect 531222 298868 531228 298920
rect 531280 298908 531286 298920
rect 536285 298911 536343 298917
rect 536285 298908 536297 298911
rect 531280 298880 536297 298908
rect 531280 298868 531286 298880
rect 536285 298877 536297 298880
rect 536331 298877 536343 298911
rect 536285 298871 536343 298877
rect 538122 298868 538128 298920
rect 538180 298908 538186 298920
rect 551554 298908 551560 298920
rect 538180 298880 551560 298908
rect 538180 298868 538186 298880
rect 551554 298868 551560 298880
rect 551612 298868 551618 298920
rect 557442 298868 557448 298920
rect 557500 298908 557506 298920
rect 564526 298908 564532 298920
rect 557500 298880 564532 298908
rect 557500 298868 557506 298880
rect 564526 298868 564532 298880
rect 564584 298868 564590 298920
rect 565722 298868 565728 298920
rect 565780 298908 565786 298920
rect 570138 298908 570144 298920
rect 565780 298880 570144 298908
rect 565780 298868 565786 298880
rect 570138 298868 570144 298880
rect 570196 298868 570202 298920
rect 425020 298812 431356 298840
rect 431405 298843 431463 298849
rect 425020 298800 425026 298812
rect 431405 298809 431417 298843
rect 431451 298840 431463 298843
rect 472802 298840 472808 298852
rect 431451 298812 472808 298840
rect 431451 298809 431463 298812
rect 431405 298803 431463 298809
rect 472802 298800 472808 298812
rect 472860 298800 472866 298852
rect 475378 298800 475384 298852
rect 475436 298840 475442 298852
rect 479429 298843 479487 298849
rect 479429 298840 479441 298843
rect 475436 298812 479441 298840
rect 475436 298800 475442 298812
rect 479429 298809 479441 298812
rect 479475 298809 479487 298843
rect 479429 298803 479487 298809
rect 480162 298800 480168 298852
rect 480220 298840 480226 298852
rect 511718 298840 511724 298852
rect 480220 298812 511724 298840
rect 480220 298800 480226 298812
rect 511718 298800 511724 298812
rect 511776 298800 511782 298852
rect 513282 298800 513288 298852
rect 513340 298840 513346 298852
rect 534442 298840 534448 298852
rect 513340 298812 534448 298840
rect 513340 298800 513346 298812
rect 534442 298800 534448 298812
rect 534500 298800 534506 298852
rect 535362 298800 535368 298852
rect 535420 298840 535426 298852
rect 549898 298840 549904 298852
rect 535420 298812 549904 298840
rect 535420 298800 535426 298812
rect 549898 298800 549904 298812
rect 549956 298800 549962 298852
rect 551278 298800 551284 298852
rect 551336 298840 551342 298852
rect 560478 298840 560484 298852
rect 551336 298812 560484 298840
rect 551336 298800 551342 298812
rect 560478 298800 560484 298812
rect 560536 298800 560542 298852
rect 7558 298732 7564 298784
rect 7616 298772 7622 298784
rect 187234 298772 187240 298784
rect 7616 298744 187240 298772
rect 7616 298732 7622 298744
rect 187234 298732 187240 298744
rect 187292 298732 187298 298784
rect 214650 298732 214656 298784
rect 214708 298772 214714 298784
rect 229370 298772 229376 298784
rect 214708 298744 229376 298772
rect 214708 298732 214714 298744
rect 229370 298732 229376 298744
rect 229428 298732 229434 298784
rect 230566 298732 230572 298784
rect 230624 298772 230630 298784
rect 267550 298772 267556 298784
rect 230624 298744 267556 298772
rect 230624 298732 230630 298744
rect 267550 298732 267556 298744
rect 267608 298732 267614 298784
rect 268378 298732 268384 298784
rect 268436 298772 268442 298784
rect 365714 298772 365720 298784
rect 268436 298744 365720 298772
rect 268436 298732 268442 298744
rect 365714 298732 365720 298744
rect 365772 298732 365778 298784
rect 367738 298732 367744 298784
rect 367796 298772 367802 298784
rect 433886 298772 433892 298784
rect 367796 298744 433892 298772
rect 367796 298732 367802 298744
rect 433886 298732 433892 298744
rect 433944 298732 433950 298784
rect 435269 298775 435327 298781
rect 435269 298741 435281 298775
rect 435315 298772 435327 298775
rect 438762 298772 438768 298784
rect 435315 298744 438768 298772
rect 435315 298741 435327 298744
rect 435269 298735 435327 298741
rect 438762 298732 438768 298744
rect 438820 298732 438826 298784
rect 438857 298775 438915 298781
rect 438857 298741 438869 298775
rect 438903 298772 438915 298775
rect 481726 298772 481732 298784
rect 438903 298744 481732 298772
rect 438903 298741 438915 298744
rect 438857 298735 438915 298741
rect 481726 298732 481732 298744
rect 481784 298732 481790 298784
rect 482922 298732 482928 298784
rect 482980 298772 482986 298784
rect 513374 298772 513380 298784
rect 482980 298744 513380 298772
rect 482980 298732 482986 298744
rect 513374 298732 513380 298744
rect 513432 298732 513438 298784
rect 516042 298732 516048 298784
rect 516100 298772 516106 298784
rect 531041 298775 531099 298781
rect 531041 298772 531053 298775
rect 516100 298744 531053 298772
rect 516100 298732 516106 298744
rect 531041 298741 531053 298744
rect 531087 298741 531099 298775
rect 531041 298735 531099 298741
rect 531133 298775 531191 298781
rect 531133 298741 531145 298775
rect 531179 298772 531191 298775
rect 537754 298772 537760 298784
rect 531179 298744 537760 298772
rect 531179 298741 531191 298744
rect 531133 298735 531191 298741
rect 537754 298732 537760 298744
rect 537812 298732 537818 298784
rect 539502 298732 539508 298784
rect 539560 298772 539566 298784
rect 552290 298772 552296 298784
rect 539560 298744 552296 298772
rect 539560 298732 539566 298744
rect 552290 298732 552296 298744
rect 552348 298732 552354 298784
rect 567102 298732 567108 298784
rect 567160 298772 567166 298784
rect 571794 298772 571800 298784
rect 567160 298744 571800 298772
rect 567160 298732 567166 298744
rect 571794 298732 571800 298744
rect 571852 298732 571858 298784
rect 582742 298772 582748 298784
rect 582703 298744 582748 298772
rect 582742 298732 582748 298744
rect 582800 298732 582806 298784
rect 101398 298664 101404 298716
rect 101456 298704 101462 298716
rect 248874 298704 248880 298716
rect 101456 298676 248880 298704
rect 101456 298664 101462 298676
rect 248874 298664 248880 298676
rect 248932 298664 248938 298716
rect 251726 298664 251732 298716
rect 251784 298704 251790 298716
rect 262674 298704 262680 298716
rect 251784 298676 262680 298704
rect 251784 298664 251790 298676
rect 262674 298664 262680 298676
rect 262732 298664 262738 298716
rect 266354 298664 266360 298716
rect 266412 298704 266418 298716
rect 278866 298704 278872 298716
rect 266412 298676 278872 298704
rect 266412 298664 266418 298676
rect 278866 298664 278872 298676
rect 278924 298664 278930 298716
rect 287790 298664 287796 298716
rect 287848 298704 287854 298716
rect 315390 298704 315396 298716
rect 287848 298676 315396 298704
rect 287848 298664 287854 298676
rect 315390 298664 315396 298676
rect 315448 298664 315454 298716
rect 329098 298664 329104 298716
rect 329156 298704 329162 298716
rect 394878 298704 394884 298716
rect 329156 298676 394884 298704
rect 329156 298664 329162 298676
rect 394878 298664 394884 298676
rect 394936 298664 394942 298716
rect 396718 298664 396724 298716
rect 396776 298704 396782 298716
rect 453298 298704 453304 298716
rect 396776 298676 453304 298704
rect 396776 298664 396782 298676
rect 453298 298664 453304 298676
rect 453356 298664 453362 298716
rect 454313 298707 454371 298713
rect 454313 298673 454325 298707
rect 454359 298704 454371 298707
rect 457346 298704 457352 298716
rect 454359 298676 457352 298704
rect 454359 298673 454371 298676
rect 454313 298667 454371 298673
rect 457346 298664 457352 298676
rect 457404 298664 457410 298716
rect 460198 298664 460204 298716
rect 460256 298704 460262 298716
rect 465534 298704 465540 298716
rect 460256 298676 465540 298704
rect 460256 298664 460262 298676
rect 465534 298664 465540 298676
rect 465592 298664 465598 298716
rect 466362 298664 466368 298716
rect 466420 298704 466426 298716
rect 502058 298704 502064 298716
rect 466420 298676 502064 298704
rect 466420 298664 466426 298676
rect 502058 298664 502064 298676
rect 502116 298664 502122 298716
rect 509142 298664 509148 298716
rect 509200 298704 509206 298716
rect 532050 298704 532056 298716
rect 509200 298676 532056 298704
rect 509200 298664 509206 298676
rect 532050 298664 532056 298676
rect 532108 298664 532114 298716
rect 533706 298704 533712 298716
rect 532160 298676 533712 298704
rect 114462 298596 114468 298648
rect 114520 298636 114526 298648
rect 261018 298636 261024 298648
rect 114520 298608 261024 298636
rect 114520 298596 114526 298608
rect 261018 298596 261024 298608
rect 261076 298596 261082 298648
rect 274542 298596 274548 298648
rect 274600 298636 274606 298648
rect 284570 298636 284576 298648
rect 274600 298608 284576 298636
rect 274600 298596 274606 298608
rect 284570 298596 284576 298608
rect 284628 298596 284634 298648
rect 298830 298596 298836 298648
rect 298888 298636 298894 298648
rect 300949 298639 301007 298645
rect 300949 298636 300961 298639
rect 298888 298608 300961 298636
rect 298888 298596 298894 298608
rect 300949 298605 300961 298608
rect 300995 298605 301007 298639
rect 300949 298599 301007 298605
rect 305822 298596 305828 298648
rect 305880 298636 305886 298648
rect 310514 298636 310520 298648
rect 305880 298608 310520 298636
rect 305880 298596 305886 298608
rect 310514 298596 310520 298608
rect 310572 298596 310578 298648
rect 324958 298596 324964 298648
rect 325016 298636 325022 298648
rect 325016 298608 373994 298636
rect 325016 298596 325022 298608
rect 121362 298528 121368 298580
rect 121420 298568 121426 298580
rect 265894 298568 265900 298580
rect 121420 298540 265900 298568
rect 121420 298528 121426 298540
rect 265894 298528 265900 298540
rect 265952 298528 265958 298580
rect 278038 298528 278044 298580
rect 278096 298568 278102 298580
rect 286781 298571 286839 298577
rect 286781 298568 286793 298571
rect 278096 298540 286793 298568
rect 278096 298528 278102 298540
rect 286781 298537 286793 298540
rect 286827 298537 286839 298571
rect 286781 298531 286839 298537
rect 305638 298528 305644 298580
rect 305696 298568 305702 298580
rect 360838 298568 360844 298580
rect 305696 298540 360844 298568
rect 305696 298528 305702 298540
rect 360838 298528 360844 298540
rect 360896 298528 360902 298580
rect 373966 298568 373994 298608
rect 384298 298596 384304 298648
rect 384356 298636 384362 298648
rect 387610 298636 387616 298648
rect 384356 298608 387616 298636
rect 384356 298596 384362 298608
rect 387610 298596 387616 298608
rect 387668 298596 387674 298648
rect 391198 298596 391204 298648
rect 391256 298636 391262 298648
rect 392486 298636 392492 298648
rect 391256 298608 392492 298636
rect 391256 298596 391262 298608
rect 392486 298596 392492 298608
rect 392544 298596 392550 298648
rect 392578 298596 392584 298648
rect 392636 298636 392642 298648
rect 397362 298636 397368 298648
rect 392636 298608 397368 298636
rect 392636 298596 392642 298608
rect 397362 298596 397368 298608
rect 397420 298596 397426 298648
rect 402238 298596 402244 298648
rect 402296 298636 402302 298648
rect 458174 298636 458180 298648
rect 402296 298608 458180 298636
rect 402296 298596 402302 298608
rect 458174 298596 458180 298608
rect 458232 298596 458238 298648
rect 482278 298596 482284 298648
rect 482336 298636 482342 298648
rect 507670 298636 507676 298648
rect 482336 298608 507676 298636
rect 482336 298596 482342 298608
rect 507670 298596 507676 298608
rect 507728 298596 507734 298648
rect 511902 298596 511908 298648
rect 511960 298636 511966 298648
rect 532160 298636 532188 298676
rect 533706 298664 533712 298676
rect 533764 298664 533770 298716
rect 538858 298664 538864 298716
rect 538916 298704 538922 298716
rect 548242 298704 548248 298716
rect 538916 298676 548248 298704
rect 538916 298664 538922 298676
rect 548242 298664 548248 298676
rect 548300 298664 548306 298716
rect 549162 298664 549168 298716
rect 549220 298704 549226 298716
rect 558822 298704 558828 298716
rect 549220 298676 558828 298704
rect 549220 298664 549226 298676
rect 558822 298664 558828 298676
rect 558880 298664 558886 298716
rect 569310 298664 569316 298716
rect 569368 298704 569374 298716
rect 570966 298704 570972 298716
rect 569368 298676 570972 298704
rect 569368 298664 569374 298676
rect 570966 298664 570972 298676
rect 571024 298664 571030 298716
rect 511960 298608 532188 298636
rect 511960 298596 511966 298608
rect 533338 298596 533344 298648
rect 533396 298636 533402 298648
rect 540974 298636 540980 298648
rect 533396 298608 540980 298636
rect 533396 298596 533402 298608
rect 540974 298596 540980 298608
rect 541032 298596 541038 298648
rect 543090 298596 543096 298648
rect 543148 298636 543154 298648
rect 553118 298636 553124 298648
rect 543148 298608 553124 298636
rect 543148 298596 543154 298608
rect 553118 298596 553124 298608
rect 553176 298596 553182 298648
rect 390002 298568 390008 298580
rect 373966 298540 390008 298568
rect 390002 298528 390008 298540
rect 390060 298528 390066 298580
rect 442169 298571 442227 298577
rect 393286 298540 442120 298568
rect 87598 298460 87604 298512
rect 87656 298500 87662 298512
rect 226978 298500 226984 298512
rect 87656 298472 226984 298500
rect 87656 298460 87662 298472
rect 226978 298460 226984 298472
rect 227036 298460 227042 298512
rect 250530 298460 250536 298512
rect 250588 298500 250594 298512
rect 253937 298503 253995 298509
rect 253937 298500 253949 298503
rect 250588 298472 253949 298500
rect 250588 298460 250594 298472
rect 253937 298469 253949 298472
rect 253983 298469 253995 298503
rect 253937 298463 253995 298469
rect 258810 298460 258816 298512
rect 258868 298500 258874 298512
rect 265161 298503 265219 298509
rect 265161 298500 265173 298503
rect 258868 298472 265173 298500
rect 258868 298460 258874 298472
rect 265161 298469 265173 298472
rect 265207 298469 265219 298503
rect 265161 298463 265219 298469
rect 338758 298460 338764 298512
rect 338816 298500 338822 298512
rect 385218 298500 385224 298512
rect 338816 298472 385224 298500
rect 338816 298460 338822 298472
rect 385218 298460 385224 298472
rect 385276 298460 385282 298512
rect 386322 298460 386328 298512
rect 386380 298500 386386 298512
rect 393286 298500 393314 298540
rect 386380 298472 393314 298500
rect 386380 298460 386386 298472
rect 396810 298460 396816 298512
rect 396868 298500 396874 298512
rect 441893 298503 441951 298509
rect 441893 298500 441905 298503
rect 396868 298472 441905 298500
rect 396868 298460 396874 298472
rect 441893 298469 441905 298472
rect 441939 298469 441951 298503
rect 441893 298463 441951 298469
rect 83458 298392 83464 298444
rect 83516 298432 83522 298444
rect 222102 298432 222108 298444
rect 83516 298404 222108 298432
rect 83516 298392 83522 298404
rect 222102 298392 222108 298404
rect 222160 298392 222166 298444
rect 317414 298392 317420 298444
rect 317472 298432 317478 298444
rect 341334 298432 341340 298444
rect 317472 298404 341340 298432
rect 317472 298392 317478 298404
rect 341334 298392 341340 298404
rect 341392 298392 341398 298444
rect 345658 298392 345664 298444
rect 345716 298432 345722 298444
rect 351181 298435 351239 298441
rect 351181 298432 351193 298435
rect 345716 298404 351193 298432
rect 345716 298392 345722 298404
rect 351181 298401 351193 298404
rect 351227 298401 351239 298435
rect 351181 298395 351239 298401
rect 358722 298392 358728 298444
rect 358780 298432 358786 298444
rect 363325 298435 363383 298441
rect 363325 298432 363337 298435
rect 358780 298404 363337 298432
rect 358780 298392 358786 298404
rect 363325 298401 363337 298404
rect 363371 298401 363383 298435
rect 363325 298395 363383 298401
rect 387702 298392 387708 298444
rect 387760 298432 387766 298444
rect 441985 298435 442043 298441
rect 441985 298432 441997 298435
rect 387760 298404 441997 298432
rect 387760 298392 387766 298404
rect 441985 298401 441997 298404
rect 442031 298401 442043 298435
rect 442092 298432 442120 298540
rect 442169 298537 442181 298571
rect 442215 298568 442227 298571
rect 443270 298568 443276 298580
rect 442215 298540 443276 298568
rect 442215 298537 442227 298540
rect 442169 298531 442227 298537
rect 443270 298528 443276 298540
rect 443328 298528 443334 298580
rect 444282 298528 444288 298580
rect 444340 298568 444346 298580
rect 450265 298571 450323 298577
rect 450265 298568 450277 298571
rect 444340 298540 450277 298568
rect 444340 298528 444346 298540
rect 450265 298537 450277 298540
rect 450311 298537 450323 298571
rect 450265 298531 450323 298537
rect 451182 298528 451188 298580
rect 451240 298568 451246 298580
rect 492306 298568 492312 298580
rect 451240 298540 492312 298568
rect 451240 298528 451246 298540
rect 492306 298528 492312 298540
rect 492364 298528 492370 298580
rect 499574 298568 499580 298580
rect 492416 298540 499580 298568
rect 442261 298503 442319 298509
rect 442261 298469 442273 298503
rect 442307 298500 442319 298503
rect 452562 298500 452568 298512
rect 442307 298472 452568 298500
rect 442307 298469 442319 298472
rect 442261 298463 442319 298469
rect 452562 298460 452568 298472
rect 452620 298460 452626 298512
rect 458082 298460 458088 298512
rect 458140 298500 458146 298512
rect 460753 298503 460811 298509
rect 460753 298500 460765 298503
rect 458140 298472 460765 298500
rect 458140 298460 458146 298472
rect 460753 298469 460765 298472
rect 460799 298469 460811 298503
rect 460753 298463 460811 298469
rect 465718 298460 465724 298512
rect 465776 298500 465782 298512
rect 489454 298500 489460 298512
rect 465776 298472 489460 298500
rect 465776 298460 465782 298472
rect 489454 298460 489460 298472
rect 489512 298460 489518 298512
rect 489886 298472 491248 298500
rect 447686 298432 447692 298444
rect 442092 298404 447692 298432
rect 441985 298395 442043 298401
rect 447686 298392 447692 298404
rect 447744 298392 447750 298444
rect 474090 298392 474096 298444
rect 474148 298432 474154 298444
rect 484210 298432 484216 298444
rect 474148 298404 484216 298432
rect 474148 298392 474154 298404
rect 484210 298392 484216 298404
rect 484268 298392 484274 298444
rect 487798 298392 487804 298444
rect 487856 298432 487862 298444
rect 489886 298432 489914 298472
rect 487856 298404 489914 298432
rect 491220 298432 491248 298472
rect 491938 298460 491944 298512
rect 491996 298500 492002 298512
rect 492416 298500 492444 298540
rect 499574 298528 499580 298540
rect 499632 298528 499638 298580
rect 502978 298528 502984 298580
rect 503036 298568 503042 298580
rect 503036 298540 521516 298568
rect 503036 298528 503042 298540
rect 491996 298472 492444 298500
rect 491996 298460 492002 298472
rect 497458 298460 497464 298512
rect 497516 298500 497522 298512
rect 510154 298500 510160 298512
rect 497516 298472 510160 298500
rect 497516 298460 497522 298472
rect 510154 298460 510160 298472
rect 510212 298460 510218 298512
rect 521488 298500 521516 298540
rect 521562 298528 521568 298580
rect 521620 298568 521626 298580
rect 528097 298571 528155 298577
rect 528097 298568 528109 298571
rect 521620 298540 528109 298568
rect 521620 298528 521626 298540
rect 528097 298537 528109 298540
rect 528143 298537 528155 298571
rect 528097 298531 528155 298537
rect 529198 298528 529204 298580
rect 529256 298568 529262 298580
rect 542630 298568 542636 298580
rect 529256 298540 542636 298568
rect 529256 298528 529262 298540
rect 542630 298528 542636 298540
rect 542688 298528 542694 298580
rect 558822 298528 558828 298580
rect 558880 298568 558886 298580
rect 566090 298568 566096 298580
rect 558880 298540 566096 298568
rect 558880 298528 558886 298540
rect 566090 298528 566096 298540
rect 566148 298528 566154 298580
rect 525518 298500 525524 298512
rect 521488 298472 525524 298500
rect 525518 298460 525524 298472
rect 525576 298460 525582 298512
rect 531041 298503 531099 298509
rect 531041 298469 531053 298503
rect 531087 298500 531099 298503
rect 536926 298500 536932 298512
rect 531087 298472 536932 298500
rect 531087 298469 531099 298472
rect 531041 298463 531099 298469
rect 536926 298460 536932 298472
rect 536984 298460 536990 298512
rect 537478 298460 537484 298512
rect 537536 298500 537542 298512
rect 545850 298500 545856 298512
rect 537536 298472 545856 298500
rect 537536 298460 537542 298472
rect 545850 298460 545856 298472
rect 545908 298460 545914 298512
rect 500773 298435 500831 298441
rect 500773 298432 500785 298435
rect 491220 298404 500785 298432
rect 487856 298392 487862 298404
rect 500773 298401 500785 298404
rect 500819 298401 500831 298435
rect 500773 298395 500831 298401
rect 500862 298392 500868 298444
rect 500920 298432 500926 298444
rect 507029 298435 507087 298441
rect 507029 298432 507041 298435
rect 500920 298404 507041 298432
rect 500920 298392 500926 298404
rect 507029 298401 507041 298404
rect 507075 298401 507087 298435
rect 507029 298395 507087 298401
rect 508498 298392 508504 298444
rect 508556 298432 508562 298444
rect 514202 298432 514208 298444
rect 508556 298404 514208 298432
rect 508556 298392 508562 298404
rect 514202 298392 514208 298404
rect 514260 298392 514266 298444
rect 520182 298392 520188 298444
rect 520240 298432 520246 298444
rect 524049 298435 524107 298441
rect 524049 298432 524061 298435
rect 520240 298404 524061 298432
rect 520240 298392 520246 298404
rect 524049 298401 524061 298404
rect 524095 298401 524107 298435
rect 524049 298395 524107 298401
rect 525058 298392 525064 298444
rect 525116 298432 525122 298444
rect 532878 298432 532884 298444
rect 525116 298404 532884 298432
rect 525116 298392 525122 298404
rect 532878 298392 532884 298404
rect 532936 298392 532942 298444
rect 536098 298392 536104 298444
rect 536156 298432 536162 298444
rect 544654 298432 544660 298444
rect 536156 298404 544660 298432
rect 536156 298392 536162 298404
rect 544654 298392 544660 298404
rect 544712 298392 544718 298444
rect 79318 298324 79324 298376
rect 79376 298364 79382 298376
rect 217226 298364 217232 298376
rect 79376 298336 217232 298364
rect 79376 298324 79382 298336
rect 217226 298324 217232 298336
rect 217284 298324 217290 298376
rect 221458 298324 221464 298376
rect 221516 298364 221522 298376
rect 224681 298367 224739 298373
rect 224681 298364 224693 298367
rect 221516 298336 224693 298364
rect 221516 298324 221522 298336
rect 224681 298333 224693 298336
rect 224727 298333 224739 298367
rect 224681 298327 224739 298333
rect 288618 298324 288624 298376
rect 288676 298364 288682 298376
rect 291010 298364 291016 298376
rect 288676 298336 291016 298364
rect 288676 298324 288682 298336
rect 291010 298324 291016 298336
rect 291068 298324 291074 298376
rect 338022 298324 338028 298376
rect 338080 298364 338086 298376
rect 340325 298367 340383 298373
rect 340325 298364 340337 298367
rect 338080 298336 340337 298364
rect 338080 298324 338086 298336
rect 340325 298333 340337 298336
rect 340371 298333 340383 298367
rect 340325 298327 340383 298333
rect 400122 298324 400128 298376
rect 400180 298364 400186 298376
rect 402333 298367 402391 298373
rect 402333 298364 402345 298367
rect 400180 298336 402345 298364
rect 400180 298324 400186 298336
rect 402333 298333 402345 298336
rect 402379 298333 402391 298367
rect 402333 298327 402391 298333
rect 411898 298324 411904 298376
rect 411956 298364 411962 298376
rect 462222 298364 462228 298376
rect 411956 298336 462228 298364
rect 411956 298324 411962 298336
rect 462222 298324 462228 298336
rect 462280 298324 462286 298376
rect 483658 298324 483664 298376
rect 483716 298364 483722 298376
rect 491113 298367 491171 298373
rect 491113 298364 491125 298367
rect 483716 298336 491125 298364
rect 483716 298324 483722 298336
rect 491113 298333 491125 298336
rect 491159 298333 491171 298367
rect 491113 298327 491171 298333
rect 491202 298324 491208 298376
rect 491260 298364 491266 298376
rect 496449 298367 496507 298373
rect 496449 298364 496461 298367
rect 491260 298336 496461 298364
rect 491260 298324 491266 298336
rect 496449 298333 496461 298336
rect 496495 298333 496507 298367
rect 496449 298327 496507 298333
rect 496722 298324 496728 298376
rect 496780 298364 496786 298376
rect 501509 298367 501567 298373
rect 501509 298364 501521 298367
rect 496780 298336 501521 298364
rect 496780 298324 496786 298336
rect 501509 298333 501521 298336
rect 501555 298333 501567 298367
rect 501509 298327 501567 298333
rect 501598 298324 501604 298376
rect 501656 298364 501662 298376
rect 510982 298364 510988 298376
rect 501656 298336 510988 298364
rect 501656 298324 501662 298336
rect 510982 298324 510988 298336
rect 511040 298324 511046 298376
rect 98638 298256 98644 298308
rect 98696 298296 98702 298308
rect 231854 298296 231860 298308
rect 98696 298268 231860 298296
rect 98696 298256 98702 298268
rect 231854 298256 231860 298268
rect 231912 298256 231918 298308
rect 416038 298256 416044 298308
rect 416096 298296 416102 298308
rect 421561 298299 421619 298305
rect 421561 298296 421573 298299
rect 416096 298268 421573 298296
rect 416096 298256 416102 298268
rect 421561 298265 421573 298268
rect 421607 298265 421619 298299
rect 421561 298259 421619 298265
rect 424318 298256 424324 298308
rect 424376 298296 424382 298308
rect 471974 298296 471980 298308
rect 424376 298268 471980 298296
rect 424376 298256 424382 298268
rect 471974 298256 471980 298268
rect 472032 298256 472038 298308
rect 480898 298256 480904 298308
rect 480956 298296 480962 298308
rect 494698 298296 494704 298308
rect 480956 298268 494704 298296
rect 480956 298256 480962 298268
rect 494698 298256 494704 298268
rect 494756 298256 494762 298308
rect 500218 298256 500224 298308
rect 500276 298296 500282 298308
rect 509326 298296 509332 298308
rect 500276 298268 509332 298296
rect 500276 298256 500282 298268
rect 509326 298256 509332 298268
rect 509384 298256 509390 298308
rect 511258 298256 511264 298308
rect 511316 298296 511322 298308
rect 529566 298296 529572 298308
rect 511316 298268 529572 298296
rect 511316 298256 511322 298268
rect 529566 298256 529572 298268
rect 529624 298256 529630 298308
rect 561582 298256 561588 298308
rect 561640 298296 561646 298308
rect 567746 298296 567752 298308
rect 561640 298268 567752 298296
rect 561640 298256 561646 298268
rect 567746 298256 567752 298268
rect 567804 298256 567810 298308
rect 105538 298188 105544 298240
rect 105596 298228 105602 298240
rect 236730 298228 236736 298240
rect 105596 298200 236736 298228
rect 105596 298188 105602 298200
rect 236730 298188 236736 298200
rect 236788 298188 236794 298240
rect 406378 298188 406384 298240
rect 406436 298228 406442 298240
rect 407114 298228 407120 298240
rect 406436 298200 407120 298228
rect 406436 298188 406442 298200
rect 407114 298188 407120 298200
rect 407172 298188 407178 298240
rect 423582 298188 423588 298240
rect 423640 298228 423646 298240
rect 431405 298231 431463 298237
rect 431405 298228 431417 298231
rect 423640 298200 431417 298228
rect 423640 298188 423646 298200
rect 431405 298197 431417 298200
rect 431451 298197 431463 298231
rect 431405 298191 431463 298197
rect 436002 298188 436008 298240
rect 436060 298228 436066 298240
rect 438857 298231 438915 298237
rect 438857 298228 438869 298231
rect 436060 298200 438869 298228
rect 436060 298188 436066 298200
rect 438857 298197 438869 298200
rect 438903 298197 438915 298231
rect 438857 298191 438915 298197
rect 447042 298188 447048 298240
rect 447100 298228 447106 298240
rect 488994 298228 489000 298240
rect 447100 298200 489000 298228
rect 447100 298188 447106 298200
rect 488994 298188 489000 298200
rect 489052 298188 489058 298240
rect 498746 298228 498752 298240
rect 489886 298200 498752 298228
rect 233878 298120 233884 298172
rect 233936 298160 233942 298172
rect 234522 298160 234528 298172
rect 233936 298132 234528 298160
rect 233936 298120 233942 298132
rect 234522 298120 234528 298132
rect 234580 298120 234586 298172
rect 263042 298120 263048 298172
rect 263100 298160 263106 298172
rect 269114 298160 269120 298172
rect 263100 298132 269120 298160
rect 263100 298120 263106 298132
rect 269114 298120 269120 298132
rect 269172 298120 269178 298172
rect 441985 298163 442043 298169
rect 441985 298129 441997 298163
rect 442031 298160 442043 298163
rect 448422 298160 448428 298172
rect 442031 298132 448428 298160
rect 442031 298129 442043 298132
rect 441985 298123 442043 298129
rect 448422 298120 448428 298132
rect 448480 298120 448486 298172
rect 479518 298120 479524 298172
rect 479576 298160 479582 298172
rect 480070 298160 480076 298172
rect 479576 298132 480076 298160
rect 479576 298120 479582 298132
rect 480070 298120 480076 298132
rect 480128 298120 480134 298172
rect 486418 298120 486424 298172
rect 486476 298160 486482 298172
rect 489886 298160 489914 298200
rect 498746 298188 498752 298200
rect 498804 298188 498810 298240
rect 504450 298228 504456 298240
rect 500236 298200 504456 298228
rect 486476 298132 489914 298160
rect 486476 298120 486482 298132
rect 492030 298120 492036 298172
rect 492088 298160 492094 298172
rect 500236 298160 500264 298200
rect 504450 298188 504456 298200
rect 504508 298188 504514 298240
rect 522298 298188 522304 298240
rect 522356 298228 522362 298240
rect 528830 298228 528836 298240
rect 522356 298200 528836 298228
rect 522356 298188 522362 298200
rect 528830 298188 528836 298200
rect 528888 298188 528894 298240
rect 565078 298188 565084 298240
rect 565136 298228 565142 298240
rect 569402 298228 569408 298240
rect 565136 298200 569408 298228
rect 565136 298188 565142 298200
rect 569402 298188 569408 298200
rect 569460 298188 569466 298240
rect 575382 298188 575388 298240
rect 575440 298228 575446 298240
rect 577498 298228 577504 298240
rect 575440 298200 577504 298228
rect 575440 298188 575446 298200
rect 577498 298188 577504 298200
rect 577556 298188 577562 298240
rect 492088 298132 500264 298160
rect 500773 298163 500831 298169
rect 492088 298120 492094 298132
rect 500773 298129 500785 298163
rect 500819 298160 500831 298163
rect 508222 298160 508228 298172
rect 500819 298132 508228 298160
rect 500819 298129 500831 298132
rect 500773 298123 500831 298129
rect 508222 298120 508228 298132
rect 508280 298120 508286 298172
rect 518158 298120 518164 298172
rect 518216 298160 518222 298172
rect 520642 298160 520648 298172
rect 518216 298132 520648 298160
rect 518216 298120 518222 298132
rect 520642 298120 520648 298132
rect 520700 298120 520706 298172
rect 554038 298120 554044 298172
rect 554096 298160 554102 298172
rect 559650 298160 559656 298172
rect 554096 298132 559656 298160
rect 554096 298120 554102 298132
rect 559650 298120 559656 298132
rect 559708 298120 559714 298172
rect 566458 298120 566464 298172
rect 566516 298160 566522 298172
rect 568574 298160 568580 298172
rect 566516 298132 568580 298160
rect 566516 298120 566522 298132
rect 568574 298120 568580 298132
rect 568632 298120 568638 298172
rect 576762 298120 576768 298172
rect 576820 298160 576826 298172
rect 578326 298160 578332 298172
rect 576820 298132 578332 298160
rect 576820 298120 576826 298132
rect 578326 298120 578332 298132
rect 578384 298120 578390 298172
rect 140682 298052 140688 298104
rect 140740 298092 140746 298104
rect 266354 298092 266360 298104
rect 140740 298064 266360 298092
rect 140740 298052 140746 298064
rect 266354 298052 266360 298064
rect 266412 298052 266418 298104
rect 341518 298052 341524 298104
rect 341576 298092 341582 298104
rect 408678 298092 408684 298104
rect 341576 298064 408684 298092
rect 341576 298052 341582 298064
rect 408678 298052 408684 298064
rect 408736 298052 408742 298104
rect 413278 298052 413284 298104
rect 413336 298092 413342 298104
rect 463878 298092 463884 298104
rect 413336 298064 463884 298092
rect 413336 298052 413342 298064
rect 463878 298052 463884 298064
rect 463936 298052 463942 298104
rect 135162 297984 135168 298036
rect 135220 298024 135226 298036
rect 263686 298024 263692 298036
rect 135220 297996 263692 298024
rect 135220 297984 135226 297996
rect 263686 297984 263692 297996
rect 263744 297984 263750 298036
rect 266998 297984 267004 298036
rect 267056 298024 267062 298036
rect 330018 298024 330024 298036
rect 267056 297996 330024 298024
rect 267056 297984 267062 297996
rect 330018 297984 330024 297996
rect 330076 297984 330082 298036
rect 343542 297984 343548 298036
rect 343600 298024 343606 298036
rect 418430 298024 418436 298036
rect 343600 297996 418436 298024
rect 343600 297984 343606 297996
rect 418430 297984 418436 297996
rect 418488 297984 418494 298036
rect 418798 297984 418804 298036
rect 418856 298024 418862 298036
rect 468754 298024 468760 298036
rect 418856 297996 468760 298024
rect 418856 297984 418862 297996
rect 468754 297984 468760 297996
rect 468812 297984 468818 298036
rect 133782 297916 133788 297968
rect 133840 297956 133846 297968
rect 273990 297956 273996 297968
rect 133840 297928 273996 297956
rect 133840 297916 133846 297928
rect 273990 297916 273996 297928
rect 274048 297916 274054 297968
rect 323578 297916 323584 297968
rect 323636 297956 323642 297968
rect 403802 297956 403808 297968
rect 323636 297928 403808 297956
rect 323636 297916 323642 297928
rect 403802 297916 403808 297928
rect 403860 297916 403866 297968
rect 407022 297916 407028 297968
rect 407080 297956 407086 297968
rect 461486 297956 461492 297968
rect 407080 297928 461492 297956
rect 407080 297916 407086 297928
rect 461486 297916 461492 297928
rect 461544 297916 461550 297968
rect 489178 297916 489184 297968
rect 489236 297956 489242 297968
rect 517054 297956 517060 297968
rect 489236 297928 517060 297956
rect 489236 297916 489242 297928
rect 517054 297916 517060 297928
rect 517112 297916 517118 297968
rect 129642 297848 129648 297900
rect 129700 297888 129706 297900
rect 271598 297888 271604 297900
rect 129700 297860 271604 297888
rect 129700 297848 129706 297860
rect 271598 297848 271604 297860
rect 271656 297848 271662 297900
rect 305730 297848 305736 297900
rect 305788 297888 305794 297900
rect 391658 297888 391664 297900
rect 305788 297860 391664 297888
rect 305788 297848 305794 297860
rect 391658 297848 391664 297860
rect 391716 297848 391722 297900
rect 401410 297888 401416 297900
rect 393286 297860 401416 297888
rect 111058 297780 111064 297832
rect 111116 297820 111122 297832
rect 257798 297820 257804 297832
rect 111116 297792 257804 297820
rect 111116 297780 111122 297792
rect 257798 297780 257804 297792
rect 257856 297780 257862 297832
rect 260098 297780 260104 297832
rect 260156 297820 260162 297832
rect 349430 297820 349436 297832
rect 260156 297792 349436 297820
rect 260156 297780 260162 297792
rect 349430 297780 349436 297792
rect 349488 297780 349494 297832
rect 360838 297780 360844 297832
rect 360896 297820 360902 297832
rect 393286 297820 393314 297860
rect 401410 297848 401416 297860
rect 401468 297848 401474 297900
rect 403618 297848 403624 297900
rect 403676 297888 403682 297900
rect 459002 297888 459008 297900
rect 403676 297860 459008 297888
rect 403676 297848 403682 297860
rect 459002 297848 459008 297860
rect 459060 297848 459066 297900
rect 461578 297848 461584 297900
rect 461636 297888 461642 297900
rect 490650 297888 490656 297900
rect 461636 297860 490656 297888
rect 461636 297848 461642 297860
rect 490650 297848 490656 297860
rect 490708 297848 490714 297900
rect 360896 297792 393314 297820
rect 360896 297780 360902 297792
rect 400858 297780 400864 297832
rect 400916 297820 400922 297832
rect 456610 297820 456616 297832
rect 400916 297792 456616 297820
rect 400916 297780 400922 297792
rect 456610 297780 456616 297792
rect 456668 297780 456674 297832
rect 468478 297780 468484 297832
rect 468536 297820 468542 297832
rect 502794 297820 502800 297832
rect 468536 297792 502800 297820
rect 468536 297780 468542 297792
rect 502794 297780 502800 297792
rect 502852 297780 502858 297832
rect 104158 297712 104164 297764
rect 104216 297752 104222 297764
rect 252922 297752 252928 297764
rect 104216 297724 252928 297752
rect 104216 297712 104222 297724
rect 252922 297712 252928 297724
rect 252980 297712 252986 297764
rect 280798 297712 280804 297764
rect 280856 297752 280862 297764
rect 373810 297752 373816 297764
rect 280856 297724 373816 297752
rect 280856 297712 280862 297724
rect 373810 297712 373816 297724
rect 373868 297712 373874 297764
rect 395982 297712 395988 297764
rect 396040 297752 396046 297764
rect 454126 297752 454132 297764
rect 396040 297724 454132 297752
rect 396040 297712 396046 297724
rect 454126 297712 454132 297724
rect 454184 297712 454190 297764
rect 471238 297712 471244 297764
rect 471296 297752 471302 297764
rect 505278 297752 505284 297764
rect 471296 297724 505284 297752
rect 471296 297712 471302 297724
rect 505278 297712 505284 297724
rect 505336 297712 505342 297764
rect 93118 297644 93124 297696
rect 93176 297684 93182 297696
rect 245654 297684 245660 297696
rect 93176 297656 245660 297684
rect 93176 297644 93182 297656
rect 245654 297644 245660 297656
rect 245712 297644 245718 297696
rect 268470 297644 268476 297696
rect 268528 297684 268534 297696
rect 361666 297684 361672 297696
rect 268528 297656 361672 297684
rect 268528 297644 268534 297656
rect 361666 297644 361672 297656
rect 361724 297644 361730 297696
rect 392670 297644 392676 297696
rect 392728 297684 392734 297696
rect 451734 297684 451740 297696
rect 392728 297656 451740 297684
rect 392728 297644 392734 297656
rect 451734 297644 451740 297656
rect 451792 297644 451798 297696
rect 464338 297644 464344 297696
rect 464396 297684 464402 297696
rect 500402 297684 500408 297696
rect 464396 297656 500408 297684
rect 464396 297644 464402 297656
rect 500402 297644 500408 297656
rect 500460 297644 500466 297696
rect 88978 297576 88984 297628
rect 89036 297616 89042 297628
rect 243170 297616 243176 297628
rect 89036 297588 243176 297616
rect 89036 297576 89042 297588
rect 243170 297576 243176 297588
rect 243228 297576 243234 297628
rect 269758 297576 269764 297628
rect 269816 297616 269822 297628
rect 366542 297616 366548 297628
rect 269816 297588 366548 297616
rect 269816 297576 269822 297588
rect 366542 297576 366548 297588
rect 366600 297576 366606 297628
rect 389818 297576 389824 297628
rect 389876 297616 389882 297628
rect 449250 297616 449256 297628
rect 389876 297588 449256 297616
rect 389876 297576 389882 297588
rect 449250 297576 449256 297588
rect 449308 297576 449314 297628
rect 457438 297576 457444 297628
rect 457496 297616 457502 297628
rect 495526 297616 495532 297628
rect 457496 297588 495532 297616
rect 457496 297576 457502 297588
rect 495526 297576 495532 297588
rect 495584 297576 495590 297628
rect 86218 297508 86224 297560
rect 86276 297548 86282 297560
rect 240778 297548 240784 297560
rect 86276 297520 240784 297548
rect 86276 297508 86282 297520
rect 240778 297508 240784 297520
rect 240836 297508 240842 297560
rect 271782 297508 271788 297560
rect 271840 297548 271846 297560
rect 368934 297548 368940 297560
rect 271840 297520 368940 297548
rect 271840 297508 271846 297520
rect 368934 297508 368940 297520
rect 368992 297508 368998 297560
rect 382182 297508 382188 297560
rect 382240 297548 382246 297560
rect 444374 297548 444380 297560
rect 382240 297520 444380 297548
rect 382240 297508 382246 297520
rect 444374 297508 444380 297520
rect 444432 297508 444438 297560
rect 453298 297508 453304 297560
rect 453356 297548 453362 297560
rect 493134 297548 493140 297560
rect 453356 297520 493140 297548
rect 453356 297508 453362 297520
rect 493134 297508 493140 297520
rect 493192 297508 493198 297560
rect 495342 297508 495348 297560
rect 495400 297548 495406 297560
rect 522022 297548 522028 297560
rect 495400 297520 522028 297548
rect 495400 297508 495406 297520
rect 522022 297508 522028 297520
rect 522080 297508 522086 297560
rect 57238 297440 57244 297492
rect 57296 297480 57302 297492
rect 211522 297480 211528 297492
rect 57296 297452 211528 297480
rect 57296 297440 57302 297452
rect 211522 297440 211528 297452
rect 211580 297440 211586 297492
rect 244918 297440 244924 297492
rect 244976 297480 244982 297492
rect 346670 297480 346676 297492
rect 244976 297452 346676 297480
rect 244976 297440 244982 297452
rect 346670 297440 346676 297452
rect 346728 297440 346734 297492
rect 378042 297440 378048 297492
rect 378100 297480 378106 297492
rect 441982 297480 441988 297492
rect 378100 297452 441988 297480
rect 378100 297440 378106 297452
rect 441982 297440 441988 297452
rect 442040 297440 442046 297492
rect 447778 297440 447784 297492
rect 447836 297480 447842 297492
rect 488258 297480 488264 297492
rect 447836 297452 488264 297480
rect 447836 297440 447842 297452
rect 488258 297440 488264 297452
rect 488316 297440 488322 297492
rect 491110 297440 491116 297492
rect 491168 297480 491174 297492
rect 519906 297480 519912 297492
rect 491168 297452 519912 297480
rect 491168 297440 491174 297452
rect 519906 297440 519912 297452
rect 519964 297440 519970 297492
rect 14458 297372 14464 297424
rect 14516 297412 14522 297424
rect 192110 297412 192116 297424
rect 14516 297384 192116 297412
rect 14516 297372 14522 297384
rect 192110 297372 192116 297384
rect 192168 297372 192174 297424
rect 242158 297372 242164 297424
rect 242216 297412 242222 297424
rect 344646 297412 344652 297424
rect 242216 297384 344652 297412
rect 242216 297372 242222 297384
rect 344646 297372 344652 297384
rect 344704 297372 344710 297424
rect 350350 297372 350356 297424
rect 350408 297412 350414 297424
rect 423306 297412 423312 297424
rect 350408 297384 423312 297412
rect 350408 297372 350414 297384
rect 423306 297372 423312 297384
rect 423364 297372 423370 297424
rect 425698 297372 425704 297424
rect 425756 297412 425762 297424
rect 473630 297412 473636 297424
rect 425756 297384 473636 297412
rect 425756 297372 425762 297384
rect 473630 297372 473636 297384
rect 473688 297372 473694 297424
rect 484302 297372 484308 297424
rect 484360 297412 484366 297424
rect 515030 297412 515036 297424
rect 484360 297384 515036 297412
rect 484360 297372 484366 297384
rect 515030 297372 515036 297384
rect 515088 297372 515094 297424
rect 179322 297304 179328 297356
rect 179380 297344 179386 297356
rect 305270 297344 305276 297356
rect 179380 297316 305276 297344
rect 179380 297304 179386 297316
rect 305270 297304 305276 297316
rect 305328 297304 305334 297356
rect 320818 297304 320824 297356
rect 320876 297344 320882 297356
rect 379514 297344 379520 297356
rect 320876 297316 379520 297344
rect 320876 297304 320882 297316
rect 379514 297304 379520 297316
rect 379572 297304 379578 297356
rect 414658 297304 414664 297356
rect 414716 297344 414722 297356
rect 466270 297344 466276 297356
rect 414716 297316 466276 297344
rect 414716 297304 414722 297316
rect 466270 297304 466276 297316
rect 466328 297304 466334 297356
rect 144822 297236 144828 297288
rect 144880 297276 144886 297288
rect 268838 297276 268844 297288
rect 144880 297248 268844 297276
rect 144880 297236 144886 297248
rect 268838 297236 268844 297248
rect 268896 297236 268902 297288
rect 356698 297236 356704 297288
rect 356756 297276 356762 297288
rect 411162 297276 411168 297288
rect 356756 297248 411168 297276
rect 356756 297236 356762 297248
rect 411162 297236 411168 297248
rect 411220 297236 411226 297288
rect 428458 297236 428464 297288
rect 428516 297276 428522 297288
rect 476022 297276 476028 297288
rect 428516 297248 476028 297276
rect 428516 297236 428522 297248
rect 476022 297236 476028 297248
rect 476080 297236 476086 297288
rect 142062 297168 142068 297220
rect 142120 297208 142126 297220
rect 262858 297208 262864 297220
rect 142120 297180 262864 297208
rect 142120 297168 142126 297180
rect 262858 297168 262864 297180
rect 262916 297168 262922 297220
rect 264238 297168 264244 297220
rect 264296 297208 264302 297220
rect 337286 297208 337292 297220
rect 264296 297180 337292 297208
rect 264296 297168 264302 297180
rect 337286 297168 337292 297180
rect 337344 297168 337350 297220
rect 370498 297168 370504 297220
rect 370556 297208 370562 297220
rect 406286 297208 406292 297220
rect 370556 297180 406292 297208
rect 370556 297168 370562 297180
rect 406286 297168 406292 297180
rect 406344 297168 406350 297220
rect 432598 297168 432604 297220
rect 432656 297208 432662 297220
rect 478506 297208 478512 297220
rect 432656 297180 478512 297208
rect 432656 297168 432662 297180
rect 478506 297168 478512 297180
rect 478564 297168 478570 297220
rect 246298 297100 246304 297152
rect 246356 297140 246362 297152
rect 332410 297140 332416 297152
rect 246356 297112 332416 297140
rect 246356 297100 246362 297112
rect 332410 297100 332416 297112
rect 332468 297100 332474 297152
rect 447870 297100 447876 297152
rect 447928 297140 447934 297152
rect 480622 297140 480628 297152
rect 447928 297112 480628 297140
rect 447928 297100 447934 297112
rect 480622 297100 480628 297112
rect 480680 297100 480686 297152
rect 250438 297032 250444 297084
rect 250496 297072 250502 297084
rect 322658 297072 322664 297084
rect 250496 297044 322664 297072
rect 250496 297032 250502 297044
rect 322658 297032 322664 297044
rect 322716 297032 322722 297084
rect 453390 297032 453396 297084
rect 453448 297072 453454 297084
rect 485774 297072 485780 297084
rect 453448 297044 485780 297072
rect 453448 297032 453454 297044
rect 485774 297032 485780 297044
rect 485832 297032 485838 297084
rect 258718 296964 258724 297016
rect 258776 297004 258782 297016
rect 325142 297004 325148 297016
rect 258776 296976 325148 297004
rect 258776 296964 258782 296976
rect 325142 296964 325148 296976
rect 325200 296964 325206 297016
rect 262858 296896 262864 296948
rect 262916 296936 262922 296948
rect 327534 296936 327540 296948
rect 262916 296908 327540 296936
rect 262916 296896 262922 296908
rect 327534 296896 327540 296908
rect 327592 296896 327598 296948
rect 177942 296624 177948 296676
rect 178000 296664 178006 296676
rect 303706 296664 303712 296676
rect 178000 296636 303712 296664
rect 178000 296624 178006 296636
rect 303706 296624 303712 296636
rect 303764 296624 303770 296676
rect 309778 296624 309784 296676
rect 309836 296664 309842 296676
rect 380986 296664 380992 296676
rect 309836 296636 380992 296664
rect 309836 296624 309842 296636
rect 380986 296624 380992 296636
rect 381044 296624 381050 296676
rect 158622 296556 158628 296608
rect 158680 296596 158686 296608
rect 288618 296596 288624 296608
rect 158680 296568 288624 296596
rect 158680 296556 158686 296568
rect 288618 296556 288624 296568
rect 288676 296556 288682 296608
rect 318058 296556 318064 296608
rect 318116 296596 318122 296608
rect 398926 296596 398932 296608
rect 318116 296568 398932 296596
rect 318116 296556 318122 296568
rect 398926 296556 398932 296568
rect 398984 296556 398990 296608
rect 147582 296488 147588 296540
rect 147640 296528 147646 296540
rect 281350 296528 281356 296540
rect 147640 296500 281356 296528
rect 147640 296488 147646 296500
rect 281350 296488 281356 296500
rect 281408 296488 281414 296540
rect 287698 296488 287704 296540
rect 287756 296528 287762 296540
rect 368474 296528 368480 296540
rect 287756 296500 368480 296528
rect 287756 296488 287762 296500
rect 368474 296488 368480 296500
rect 368532 296488 368538 296540
rect 151722 296420 151728 296472
rect 151780 296460 151786 296472
rect 285766 296460 285772 296472
rect 151780 296432 285772 296460
rect 151780 296420 151786 296432
rect 285766 296420 285772 296432
rect 285824 296420 285830 296472
rect 304258 296420 304264 296472
rect 304316 296460 304322 296472
rect 386506 296460 386512 296472
rect 304316 296432 386512 296460
rect 304316 296420 304322 296432
rect 386506 296420 386512 296432
rect 386564 296420 386570 296472
rect 113082 296352 113088 296404
rect 113140 296392 113146 296404
rect 259546 296392 259552 296404
rect 113140 296364 259552 296392
rect 113140 296352 113146 296364
rect 259546 296352 259552 296364
rect 259604 296352 259610 296404
rect 273898 296352 273904 296404
rect 273956 296392 273962 296404
rect 357526 296392 357532 296404
rect 273956 296364 357532 296392
rect 273956 296352 273962 296364
rect 357526 296352 357532 296364
rect 357584 296352 357590 296404
rect 108298 296284 108304 296336
rect 108356 296324 108362 296336
rect 255406 296324 255412 296336
rect 108356 296296 255412 296324
rect 108356 296284 108362 296296
rect 255406 296284 255412 296296
rect 255464 296284 255470 296336
rect 298738 296284 298744 296336
rect 298796 296324 298802 296336
rect 383654 296324 383660 296336
rect 298796 296296 383660 296324
rect 298796 296284 298802 296296
rect 383654 296284 383660 296296
rect 383712 296284 383718 296336
rect 99282 296216 99288 296268
rect 99340 296256 99346 296268
rect 249794 296256 249800 296268
rect 99340 296228 249800 296256
rect 99340 296216 99346 296228
rect 249794 296216 249800 296228
rect 249852 296216 249858 296268
rect 286318 296216 286324 296268
rect 286376 296256 286382 296268
rect 376846 296256 376852 296268
rect 286376 296228 376852 296256
rect 286376 296216 286382 296228
rect 376846 296216 376852 296228
rect 376904 296216 376910 296268
rect 95142 296148 95148 296200
rect 95200 296188 95206 296200
rect 246942 296188 246948 296200
rect 95200 296160 246948 296188
rect 95200 296148 95206 296160
rect 246942 296148 246948 296160
rect 247000 296148 247006 296200
rect 262950 296148 262956 296200
rect 263008 296188 263014 296200
rect 361574 296188 361580 296200
rect 263008 296160 361580 296188
rect 263008 296148 263014 296160
rect 361574 296148 361580 296160
rect 361632 296148 361638 296200
rect 376018 296148 376024 296200
rect 376076 296188 376082 296200
rect 432046 296188 432052 296200
rect 376076 296160 432052 296188
rect 376076 296148 376082 296160
rect 432046 296148 432052 296160
rect 432104 296148 432110 296200
rect 54478 296080 54484 296132
rect 54536 296120 54542 296132
rect 214006 296120 214012 296132
rect 54536 296092 214012 296120
rect 54536 296080 54542 296092
rect 214006 296080 214012 296092
rect 214064 296080 214070 296132
rect 240778 296080 240784 296132
rect 240836 296120 240842 296132
rect 343634 296120 343640 296132
rect 240836 296092 343640 296120
rect 240836 296080 240842 296092
rect 343634 296080 343640 296092
rect 343692 296080 343698 296132
rect 370590 296080 370596 296132
rect 370648 296120 370654 296132
rect 434806 296120 434812 296132
rect 370648 296092 434812 296120
rect 370648 296080 370654 296092
rect 434806 296080 434812 296092
rect 434864 296080 434870 296132
rect 47578 296012 47584 296064
rect 47636 296052 47642 296064
rect 208394 296052 208400 296064
rect 47636 296024 208400 296052
rect 47636 296012 47642 296024
rect 208394 296012 208400 296024
rect 208452 296012 208458 296064
rect 223482 296012 223488 296064
rect 223540 296052 223546 296064
rect 335446 296052 335452 296064
rect 223540 296024 335452 296052
rect 223540 296012 223546 296024
rect 335446 296012 335452 296024
rect 335504 296012 335510 296064
rect 375282 296012 375288 296064
rect 375340 296052 375346 296064
rect 440326 296052 440332 296064
rect 375340 296024 440332 296052
rect 375340 296012 375346 296024
rect 440326 296012 440332 296024
rect 440384 296012 440390 296064
rect 25498 295944 25504 295996
rect 25556 295984 25562 295996
rect 197446 295984 197452 295996
rect 25556 295956 197452 295984
rect 25556 295944 25562 295956
rect 197446 295944 197452 295956
rect 197504 295944 197510 295996
rect 209682 295944 209688 295996
rect 209740 295984 209746 295996
rect 325786 295984 325792 295996
rect 209740 295956 325792 295984
rect 209740 295944 209746 295956
rect 325786 295944 325792 295956
rect 325844 295944 325850 295996
rect 336642 295944 336648 295996
rect 336700 295984 336706 295996
rect 412726 295984 412732 295996
rect 336700 295956 412732 295984
rect 336700 295944 336706 295956
rect 412726 295944 412732 295956
rect 412784 295944 412790 295996
rect 439498 295944 439504 295996
rect 439556 295984 439562 295996
rect 483106 295984 483112 295996
rect 439556 295956 483112 295984
rect 439556 295944 439562 295956
rect 483106 295944 483112 295956
rect 483164 295944 483170 295996
rect 148962 295876 148968 295928
rect 149020 295916 149026 295928
rect 274542 295916 274548 295928
rect 149020 295888 274548 295916
rect 149020 295876 149026 295888
rect 274542 295876 274548 295888
rect 274600 295876 274606 295928
rect 291838 295876 291844 295928
rect 291896 295916 291902 295928
rect 371326 295916 371332 295928
rect 291896 295888 371332 295916
rect 291896 295876 291902 295888
rect 371326 295876 371332 295888
rect 371384 295876 371390 295928
rect 256050 295808 256056 295860
rect 256108 295848 256114 295860
rect 338206 295848 338212 295860
rect 256108 295820 338212 295848
rect 256108 295808 256114 295820
rect 338206 295808 338212 295820
rect 338264 295808 338270 295860
rect 251818 295740 251824 295792
rect 251876 295780 251882 295792
rect 332594 295780 332600 295792
rect 251876 295752 332600 295780
rect 251876 295740 251882 295752
rect 332594 295740 332600 295752
rect 332652 295740 332658 295792
rect 124122 294856 124128 294908
rect 124180 294896 124186 294908
rect 230566 294896 230572 294908
rect 124180 294868 230572 294896
rect 124180 294856 124186 294868
rect 230566 294856 230572 294868
rect 230624 294856 230630 294908
rect 117222 294788 117228 294840
rect 117280 294828 117286 294840
rect 251726 294828 251732 294840
rect 117280 294800 251732 294828
rect 117280 294788 117286 294800
rect 251726 294788 251732 294800
rect 251784 294788 251790 294840
rect 119982 294720 119988 294772
rect 120040 294760 120046 294772
rect 258074 294760 258080 294772
rect 120040 294732 258080 294760
rect 120040 294720 120046 294732
rect 258074 294720 258080 294732
rect 258132 294720 258138 294772
rect 51810 294652 51816 294704
rect 51868 294692 51874 294704
rect 205726 294692 205732 294704
rect 51868 294664 205732 294692
rect 51868 294652 51874 294664
rect 205726 294652 205732 294664
rect 205784 294652 205790 294704
rect 32398 294584 32404 294636
rect 32456 294624 32462 294636
rect 201586 294624 201592 294636
rect 32456 294596 201592 294624
rect 32456 294584 32462 294596
rect 201586 294584 201592 294596
rect 201644 294584 201650 294636
rect 231762 294584 231768 294636
rect 231820 294624 231826 294636
rect 317414 294624 317420 294636
rect 231820 294596 317420 294624
rect 231820 294584 231826 294596
rect 317414 294584 317420 294596
rect 317472 294584 317478 294636
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 51718 293944 51724 293956
rect 3108 293916 51724 293944
rect 3108 293904 3114 293916
rect 51718 293904 51724 293916
rect 51776 293904 51782 293956
rect 582650 258924 582656 258936
rect 582611 258896 582656 258924
rect 582650 258884 582656 258896
rect 582708 258884 582714 258936
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 40678 255252 40684 255264
rect 3200 255224 40684 255252
rect 3200 255212 3206 255224
rect 40678 255212 40684 255224
rect 40736 255212 40742 255264
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 39390 241448 39396 241460
rect 3568 241420 39396 241448
rect 3568 241408 3574 241420
rect 39390 241408 39396 241420
rect 39448 241408 39454 241460
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 137278 202824 137284 202836
rect 3108 202796 137284 202824
rect 3108 202784 3114 202796
rect 137278 202784 137284 202796
rect 137336 202784 137342 202836
rect 137922 202104 137928 202156
rect 137980 202144 137986 202156
rect 276106 202144 276112 202156
rect 137980 202116 276112 202144
rect 137980 202104 137986 202116
rect 276106 202104 276112 202116
rect 276164 202104 276170 202156
rect 276658 202104 276664 202156
rect 276716 202144 276722 202156
rect 367186 202144 367192 202156
rect 276716 202116 367192 202144
rect 276716 202104 276722 202116
rect 367186 202104 367192 202116
rect 367244 202104 367250 202156
rect 153102 188300 153108 188352
rect 153160 188340 153166 188352
rect 285674 188340 285680 188352
rect 153160 188312 285680 188340
rect 153160 188300 153166 188312
rect 285674 188300 285680 188312
rect 285732 188300 285738 188352
rect 582558 165900 582564 165912
rect 582519 165872 582564 165900
rect 582558 165860 582564 165872
rect 582616 165860 582622 165912
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 180058 164200 180064 164212
rect 3292 164172 180064 164200
rect 3292 164160 3298 164172
rect 180058 164160 180064 164172
rect 180116 164160 180122 164212
rect 582466 152708 582472 152720
rect 582427 152680 582472 152708
rect 582466 152668 582472 152680
rect 582524 152668 582530 152720
rect 274082 141380 274088 141432
rect 274140 141420 274146 141432
rect 340966 141420 340972 141432
rect 274140 141392 340972 141420
rect 274140 141380 274146 141392
rect 340966 141380 340972 141392
rect 341024 141380 341030 141432
rect 240962 140020 240968 140072
rect 241020 140060 241026 140072
rect 320266 140060 320272 140072
rect 241020 140032 320272 140060
rect 241020 140020 241026 140032
rect 320266 140020 320272 140032
rect 320324 140020 320330 140072
rect 240870 139340 240876 139392
rect 240928 139380 240934 139392
rect 579798 139380 579804 139392
rect 240928 139352 579804 139380
rect 240928 139340 240934 139352
rect 579798 139340 579804 139352
rect 579856 139340 579862 139392
rect 182910 113092 182916 113144
rect 182968 113132 182974 113144
rect 579982 113132 579988 113144
rect 182968 113104 579988 113132
rect 182968 113092 182974 113104
rect 579982 113092 579988 113104
rect 580040 113092 580046 113144
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 15838 111772 15844 111784
rect 3476 111744 15844 111772
rect 3476 111732 3482 111744
rect 15838 111732 15844 111744
rect 15896 111732 15902 111784
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 36538 97968 36544 97980
rect 3476 97940 36544 97968
rect 3476 97928 3482 97940
rect 36538 97928 36544 97940
rect 36596 97928 36602 97980
rect 183002 86912 183008 86964
rect 183060 86952 183066 86964
rect 580166 86952 580172 86964
rect 183060 86924 580172 86952
rect 183060 86912 183066 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 39298 85524 39304 85536
rect 3200 85496 39304 85524
rect 3200 85484 3206 85496
rect 39298 85484 39304 85496
rect 39356 85484 39362 85536
rect 181898 73108 181904 73160
rect 181956 73148 181962 73160
rect 580166 73148 580172 73160
rect 181956 73120 580172 73148
rect 181956 73108 181962 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 22738 71720 22744 71732
rect 3476 71692 22744 71720
rect 3476 71680 3482 71692
rect 22738 71680 22744 71692
rect 22796 71680 22802 71732
rect 155862 48968 155868 49020
rect 155920 49008 155926 49020
rect 288526 49008 288532 49020
rect 155920 48980 288532 49008
rect 155920 48968 155926 48980
rect 288526 48968 288532 48980
rect 288584 48968 288590 49020
rect 183094 46860 183100 46912
rect 183152 46900 183158 46912
rect 580166 46900 580172 46912
rect 183152 46872 580172 46900
rect 183152 46860 183158 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 61378 45540 61384 45552
rect 3476 45512 61384 45540
rect 3476 45500 3482 45512
rect 61378 45500 61384 45512
rect 61436 45500 61442 45552
rect 39298 39312 39304 39364
rect 39356 39352 39362 39364
rect 204346 39352 204352 39364
rect 39356 39324 204352 39352
rect 39356 39312 39362 39324
rect 204346 39312 204352 39324
rect 204404 39312 204410 39364
rect 181990 33056 181996 33108
rect 182048 33096 182054 33108
rect 579798 33096 579804 33108
rect 182048 33068 579804 33096
rect 182048 33056 182054 33068
rect 579798 33056 579804 33068
rect 579856 33056 579862 33108
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 583754 20652 583760 20664
rect 3476 20624 583760 20652
rect 3476 20612 3482 20624
rect 583754 20612 583760 20624
rect 583812 20612 583818 20664
rect 182082 20544 182088 20596
rect 182140 20584 182146 20596
rect 580166 20584 580172 20596
rect 182140 20556 580172 20584
rect 182140 20544 182146 20556
rect 580166 20544 580172 20556
rect 580224 20544 580230 20596
rect 22738 19932 22744 19984
rect 22796 19972 22802 19984
rect 194594 19972 194600 19984
rect 22796 19944 194600 19972
rect 22796 19932 22802 19944
rect 194594 19932 194600 19944
rect 194652 19932 194658 19984
rect 312630 18572 312636 18624
rect 312688 18612 312694 18624
rect 396166 18612 396172 18624
rect 312688 18584 396172 18612
rect 312688 18572 312694 18584
rect 396166 18572 396172 18584
rect 396224 18572 396230 18624
rect 195882 17212 195888 17264
rect 195940 17252 195946 17264
rect 316126 17252 316132 17264
rect 195940 17224 316132 17252
rect 195940 17212 195946 17224
rect 316126 17212 316132 17224
rect 316184 17212 316190 17264
rect 289078 14628 289084 14680
rect 289136 14668 289142 14680
rect 373994 14668 374000 14680
rect 289136 14640 374000 14668
rect 289136 14628 289142 14640
rect 373994 14628 374000 14640
rect 374052 14628 374058 14680
rect 271138 14560 271144 14612
rect 271196 14600 271202 14612
rect 358906 14600 358912 14612
rect 271196 14572 358912 14600
rect 271196 14560 271202 14572
rect 358906 14560 358912 14572
rect 358964 14560 358970 14612
rect 267090 14492 267096 14544
rect 267148 14532 267154 14544
rect 364334 14532 364340 14544
rect 267148 14504 364340 14532
rect 267148 14492 267154 14504
rect 364334 14492 364340 14504
rect 364392 14492 364398 14544
rect 81342 14424 81348 14476
rect 81400 14464 81406 14476
rect 237466 14464 237472 14476
rect 81400 14436 237472 14464
rect 81400 14424 81406 14436
rect 237466 14424 237472 14436
rect 237524 14424 237530 14476
rect 238018 14424 238024 14476
rect 238076 14464 238082 14476
rect 339586 14464 339592 14476
rect 238076 14436 339592 14464
rect 238076 14424 238082 14436
rect 339586 14424 339592 14436
rect 339644 14424 339650 14476
rect 169662 13132 169668 13184
rect 169720 13172 169726 13184
rect 250530 13172 250536 13184
rect 169720 13144 250536 13172
rect 169720 13132 169726 13144
rect 250530 13132 250536 13144
rect 250588 13132 250594 13184
rect 253382 13132 253388 13184
rect 253440 13172 253446 13184
rect 334066 13172 334072 13184
rect 253440 13144 334072 13172
rect 253440 13132 253446 13144
rect 334066 13132 334072 13144
rect 334124 13132 334130 13184
rect 200022 13064 200028 13116
rect 200080 13104 200086 13116
rect 312538 13104 312544 13116
rect 200080 13076 312544 13104
rect 200080 13064 200086 13076
rect 312538 13064 312544 13076
rect 312596 13064 312602 13116
rect 197262 12180 197268 12232
rect 197320 12220 197326 12232
rect 273990 12220 273996 12232
rect 197320 12192 273996 12220
rect 197320 12180 197326 12192
rect 273990 12180 273996 12192
rect 274048 12180 274054 12232
rect 251082 12112 251088 12164
rect 251140 12152 251146 12164
rect 353386 12152 353392 12164
rect 251140 12124 353392 12152
rect 251140 12112 251146 12124
rect 353386 12112 353392 12124
rect 353444 12112 353450 12164
rect 188982 12044 188988 12096
rect 189040 12084 189046 12096
rect 300118 12084 300124 12096
rect 189040 12056 300124 12084
rect 189040 12044 189046 12056
rect 300118 12044 300124 12056
rect 300176 12044 300182 12096
rect 132402 11976 132408 12028
rect 132460 12016 132466 12028
rect 253290 12016 253296 12028
rect 132460 11988 253296 12016
rect 132460 11976 132466 11988
rect 253290 11976 253296 11988
rect 253348 11976 253354 12028
rect 182082 11908 182088 11960
rect 182140 11948 182146 11960
rect 306466 11948 306472 11960
rect 182140 11920 306472 11948
rect 182140 11908 182146 11920
rect 306466 11908 306472 11920
rect 306524 11908 306530 11960
rect 176562 11840 176568 11892
rect 176620 11880 176626 11892
rect 302326 11880 302332 11892
rect 176620 11852 302332 11880
rect 176620 11840 176626 11852
rect 302326 11840 302332 11852
rect 302384 11840 302390 11892
rect 359458 11840 359464 11892
rect 359516 11880 359522 11892
rect 427906 11880 427912 11892
rect 359516 11852 427912 11880
rect 359516 11840 359522 11852
rect 427906 11840 427912 11852
rect 427964 11840 427970 11892
rect 154206 11772 154212 11824
rect 154264 11812 154270 11824
rect 288434 11812 288440 11824
rect 154264 11784 288440 11812
rect 154264 11772 154270 11784
rect 288434 11772 288440 11784
rect 288492 11772 288498 11824
rect 354582 11772 354588 11824
rect 354640 11812 354646 11824
rect 425054 11812 425060 11824
rect 354640 11784 425060 11812
rect 354640 11772 354646 11784
rect 425054 11772 425060 11784
rect 425112 11772 425118 11824
rect 144730 11704 144736 11756
rect 144788 11744 144794 11756
rect 281534 11744 281540 11756
rect 144788 11716 281540 11744
rect 144788 11704 144794 11716
rect 281534 11704 281540 11716
rect 281592 11704 281598 11756
rect 300762 11704 300768 11756
rect 300820 11744 300826 11756
rect 389266 11744 389272 11756
rect 300820 11716 389272 11744
rect 300820 11704 300826 11716
rect 389266 11704 389272 11716
rect 389324 11704 389330 11756
rect 194502 10956 194508 11008
rect 194560 10996 194566 11008
rect 287790 10996 287796 11008
rect 194560 10968 287796 10996
rect 194560 10956 194566 10968
rect 287790 10956 287796 10968
rect 287848 10956 287854 11008
rect 161290 10888 161296 10940
rect 161348 10928 161354 10940
rect 258810 10928 258816 10940
rect 161348 10900 258816 10928
rect 161348 10888 161354 10900
rect 258810 10888 258816 10900
rect 258868 10888 258874 10940
rect 259362 10888 259368 10940
rect 259420 10928 259426 10940
rect 358814 10928 358820 10940
rect 259420 10900 358820 10928
rect 259420 10888 259426 10900
rect 358814 10888 358820 10900
rect 358872 10888 358878 10940
rect 165522 10820 165528 10872
rect 165580 10860 165586 10872
rect 253198 10860 253204 10872
rect 165580 10832 253204 10860
rect 165580 10820 165586 10832
rect 253198 10820 253204 10832
rect 253256 10820 253262 10872
rect 253842 10820 253848 10872
rect 253900 10860 253906 10872
rect 356054 10860 356060 10872
rect 253900 10832 356060 10860
rect 253900 10820 253906 10832
rect 356054 10820 356060 10832
rect 356112 10820 356118 10872
rect 190362 10752 190368 10804
rect 190420 10792 190426 10804
rect 296070 10792 296076 10804
rect 190420 10764 296076 10792
rect 190420 10752 190426 10764
rect 296070 10752 296076 10764
rect 296128 10752 296134 10804
rect 183462 10684 183468 10736
rect 183520 10724 183526 10736
rect 298830 10724 298836 10736
rect 183520 10696 298836 10724
rect 183520 10684 183526 10696
rect 298830 10684 298836 10696
rect 298888 10684 298894 10736
rect 186130 10616 186136 10668
rect 186188 10656 186194 10668
rect 305822 10656 305828 10668
rect 186188 10628 305828 10656
rect 186188 10616 186194 10628
rect 305822 10616 305828 10628
rect 305880 10616 305886 10668
rect 126882 10548 126888 10600
rect 126940 10588 126946 10600
rect 263042 10588 263048 10600
rect 126940 10560 263048 10588
rect 126940 10548 126946 10560
rect 263042 10548 263048 10560
rect 263100 10548 263106 10600
rect 269850 10548 269856 10600
rect 269908 10588 269914 10600
rect 352006 10588 352012 10600
rect 269908 10560 352012 10588
rect 269908 10548 269914 10560
rect 352006 10548 352012 10560
rect 352064 10548 352070 10600
rect 136450 10480 136456 10532
rect 136508 10520 136514 10532
rect 276014 10520 276020 10532
rect 136508 10492 276020 10520
rect 136508 10480 136514 10492
rect 276014 10480 276020 10492
rect 276072 10480 276078 10532
rect 296622 10480 296628 10532
rect 296680 10520 296686 10532
rect 385126 10520 385132 10532
rect 296680 10492 385132 10520
rect 296680 10480 296686 10492
rect 385126 10480 385132 10492
rect 385184 10480 385190 10532
rect 122742 10412 122748 10464
rect 122800 10452 122806 10464
rect 266446 10452 266452 10464
rect 122800 10424 266452 10452
rect 122800 10412 122806 10424
rect 266446 10412 266452 10424
rect 266504 10412 266510 10464
rect 276750 10412 276756 10464
rect 276808 10452 276814 10464
rect 371234 10452 371240 10464
rect 276808 10424 371240 10452
rect 276808 10412 276814 10424
rect 371234 10412 371240 10424
rect 371292 10412 371298 10464
rect 119798 10344 119804 10396
rect 119856 10384 119862 10396
rect 263594 10384 263600 10396
rect 119856 10356 263600 10384
rect 119856 10344 119862 10356
rect 263594 10344 263600 10356
rect 263652 10344 263658 10396
rect 264882 10344 264888 10396
rect 264940 10384 264946 10396
rect 363046 10384 363052 10396
rect 264940 10356 363052 10384
rect 264940 10344 264946 10356
rect 363046 10344 363052 10356
rect 363104 10344 363110 10396
rect 363598 10344 363604 10396
rect 363656 10384 363662 10396
rect 430666 10384 430672 10396
rect 363656 10356 430672 10384
rect 363656 10344 363662 10356
rect 430666 10344 430672 10356
rect 430724 10344 430730 10396
rect 3418 10276 3424 10328
rect 3476 10316 3482 10328
rect 582377 10319 582435 10325
rect 582377 10316 582389 10319
rect 3476 10288 582389 10316
rect 3476 10276 3482 10288
rect 582377 10285 582389 10288
rect 582423 10285 582435 10319
rect 582377 10279 582435 10285
rect 172422 10208 172428 10260
rect 172480 10248 172486 10260
rect 246390 10248 246396 10260
rect 172480 10220 246396 10248
rect 172480 10208 172486 10220
rect 246390 10208 246396 10220
rect 246448 10208 246454 10260
rect 156598 9596 156604 9648
rect 156656 9636 156662 9648
rect 289906 9636 289912 9648
rect 156656 9608 289912 9636
rect 156656 9596 156662 9608
rect 289906 9596 289912 9608
rect 289964 9596 289970 9648
rect 149514 9528 149520 9580
rect 149572 9568 149578 9580
rect 284386 9568 284392 9580
rect 149572 9540 284392 9568
rect 149572 9528 149578 9540
rect 284386 9528 284392 9540
rect 284444 9528 284450 9580
rect 153010 9460 153016 9512
rect 153068 9500 153074 9512
rect 287054 9500 287060 9512
rect 153068 9472 287060 9500
rect 153068 9460 153074 9472
rect 287054 9460 287060 9472
rect 287112 9460 287118 9512
rect 145926 9392 145932 9444
rect 145984 9432 145990 9444
rect 283006 9432 283012 9444
rect 145984 9404 283012 9432
rect 145984 9392 145990 9404
rect 283006 9392 283012 9404
rect 283064 9392 283070 9444
rect 142430 9324 142436 9376
rect 142488 9364 142494 9376
rect 280246 9364 280252 9376
rect 142488 9336 280252 9364
rect 142488 9324 142494 9336
rect 280246 9324 280252 9336
rect 280304 9324 280310 9376
rect 138842 9256 138848 9308
rect 138900 9296 138906 9308
rect 277394 9296 277400 9308
rect 138900 9268 277400 9296
rect 138900 9256 138906 9268
rect 277394 9256 277400 9268
rect 277452 9256 277458 9308
rect 135254 9188 135260 9240
rect 135312 9228 135318 9240
rect 274726 9228 274732 9240
rect 135312 9200 274732 9228
rect 135312 9188 135318 9200
rect 274726 9188 274732 9200
rect 274784 9188 274790 9240
rect 115198 9120 115204 9172
rect 115256 9160 115262 9172
rect 260926 9160 260932 9172
rect 115256 9132 260932 9160
rect 115256 9120 115262 9132
rect 260926 9120 260932 9132
rect 260984 9120 260990 9172
rect 108114 9052 108120 9104
rect 108172 9092 108178 9104
rect 256694 9092 256700 9104
rect 108172 9064 256700 9092
rect 108172 9052 108178 9064
rect 256694 9052 256700 9064
rect 256752 9052 256758 9104
rect 111610 8984 111616 9036
rect 111668 9024 111674 9036
rect 259454 9024 259460 9036
rect 111668 8996 259460 9024
rect 111668 8984 111674 8996
rect 259454 8984 259460 8996
rect 259512 8984 259518 9036
rect 104526 8916 104532 8968
rect 104584 8956 104590 8968
rect 253934 8956 253940 8968
rect 104584 8928 253940 8956
rect 104584 8916 104590 8928
rect 253934 8916 253940 8928
rect 253992 8916 253998 8968
rect 160094 8848 160100 8900
rect 160152 8888 160158 8900
rect 292666 8888 292672 8900
rect 160152 8860 292672 8888
rect 160152 8848 160158 8860
rect 292666 8848 292672 8860
rect 292724 8848 292730 8900
rect 206186 8780 206192 8832
rect 206244 8820 206250 8832
rect 324314 8820 324320 8832
rect 206244 8792 324320 8820
rect 206244 8780 206250 8792
rect 324314 8780 324320 8792
rect 324372 8780 324378 8832
rect 213362 8712 213368 8764
rect 213420 8752 213426 8764
rect 328454 8752 328460 8764
rect 213420 8724 328460 8752
rect 213420 8712 213426 8724
rect 328454 8712 328460 8724
rect 328512 8712 328518 8764
rect 209774 8644 209780 8696
rect 209832 8684 209838 8696
rect 325694 8684 325700 8696
rect 209832 8656 325700 8684
rect 209832 8644 209838 8656
rect 325694 8644 325700 8656
rect 325752 8644 325758 8696
rect 216858 8576 216864 8628
rect 216916 8616 216922 8628
rect 331214 8616 331220 8628
rect 216916 8588 331220 8616
rect 216916 8576 216922 8588
rect 331214 8576 331220 8588
rect 331272 8576 331278 8628
rect 220446 8508 220452 8560
rect 220504 8548 220510 8560
rect 333974 8548 333980 8560
rect 220504 8520 333980 8548
rect 220504 8508 220510 8520
rect 333974 8508 333980 8520
rect 334032 8508 334038 8560
rect 227530 8440 227536 8492
rect 227588 8480 227594 8492
rect 338114 8480 338120 8492
rect 227588 8452 338120 8480
rect 227588 8440 227594 8452
rect 338114 8440 338120 8452
rect 338172 8440 338178 8492
rect 223942 8372 223948 8424
rect 224000 8412 224006 8424
rect 335354 8412 335360 8424
rect 224000 8384 335360 8412
rect 224000 8372 224006 8384
rect 335354 8372 335360 8384
rect 335412 8372 335418 8424
rect 73798 8236 73804 8288
rect 73856 8276 73862 8288
rect 233326 8276 233332 8288
rect 73856 8248 233332 8276
rect 73856 8236 73862 8248
rect 233326 8236 233332 8248
rect 233384 8236 233390 8288
rect 70302 8168 70308 8220
rect 70360 8208 70366 8220
rect 230474 8208 230480 8220
rect 70360 8180 230480 8208
rect 70360 8168 70366 8180
rect 230474 8168 230480 8180
rect 230532 8168 230538 8220
rect 66714 8100 66720 8152
rect 66772 8140 66778 8152
rect 227806 8140 227812 8152
rect 66772 8112 227812 8140
rect 66772 8100 66778 8112
rect 227806 8100 227812 8112
rect 227864 8100 227870 8152
rect 63218 8032 63224 8084
rect 63276 8072 63282 8084
rect 225046 8072 225052 8084
rect 63276 8044 225052 8072
rect 63276 8032 63282 8044
rect 225046 8032 225052 8044
rect 225104 8032 225110 8084
rect 59630 7964 59636 8016
rect 59688 8004 59694 8016
rect 223666 8004 223672 8016
rect 59688 7976 223672 8004
rect 59688 7964 59694 7976
rect 223666 7964 223672 7976
rect 223724 7964 223730 8016
rect 56042 7896 56048 7948
rect 56100 7936 56106 7948
rect 220906 7936 220912 7948
rect 56100 7908 220912 7936
rect 56100 7896 56106 7908
rect 220906 7896 220912 7908
rect 220964 7896 220970 7948
rect 251174 7896 251180 7948
rect 251232 7936 251238 7948
rect 354766 7936 354772 7948
rect 251232 7908 354772 7936
rect 251232 7896 251238 7908
rect 354766 7896 354772 7908
rect 354824 7896 354830 7948
rect 52546 7828 52552 7880
rect 52604 7868 52610 7880
rect 218146 7868 218152 7880
rect 52604 7840 218152 7868
rect 52604 7828 52610 7840
rect 218146 7828 218152 7840
rect 218204 7828 218210 7880
rect 247586 7828 247592 7880
rect 247644 7868 247650 7880
rect 351914 7868 351920 7880
rect 247644 7840 351920 7868
rect 247644 7828 247650 7840
rect 351914 7828 351920 7840
rect 351972 7828 351978 7880
rect 48958 7760 48964 7812
rect 49016 7800 49022 7812
rect 215386 7800 215392 7812
rect 49016 7772 215392 7800
rect 49016 7760 49022 7772
rect 215386 7760 215392 7772
rect 215444 7760 215450 7812
rect 244090 7760 244096 7812
rect 244148 7800 244154 7812
rect 349154 7800 349160 7812
rect 244148 7772 349160 7800
rect 244148 7760 244154 7772
rect 349154 7760 349160 7772
rect 349212 7760 349218 7812
rect 44266 7692 44272 7744
rect 44324 7732 44330 7744
rect 212534 7732 212540 7744
rect 44324 7704 212540 7732
rect 44324 7692 44330 7704
rect 212534 7692 212540 7704
rect 212592 7692 212598 7744
rect 240502 7692 240508 7744
rect 240560 7732 240566 7744
rect 347866 7732 347872 7744
rect 240560 7704 347872 7732
rect 240560 7692 240566 7704
rect 347866 7692 347872 7704
rect 347924 7692 347930 7744
rect 40678 7624 40684 7676
rect 40736 7664 40742 7676
rect 209866 7664 209872 7676
rect 40736 7636 209872 7664
rect 40736 7624 40742 7636
rect 209866 7624 209872 7636
rect 209924 7624 209930 7676
rect 233418 7624 233424 7676
rect 233476 7664 233482 7676
rect 342254 7664 342260 7676
rect 233476 7636 342260 7664
rect 233476 7624 233482 7636
rect 342254 7624 342260 7636
rect 342312 7624 342318 7676
rect 37182 7556 37188 7608
rect 37240 7596 37246 7608
rect 207106 7596 207112 7608
rect 37240 7568 207112 7596
rect 37240 7556 37246 7568
rect 207106 7556 207112 7568
rect 207164 7556 207170 7608
rect 237006 7556 237012 7608
rect 237064 7596 237070 7608
rect 345106 7596 345112 7608
rect 237064 7568 345112 7596
rect 237064 7556 237070 7568
rect 345106 7556 345112 7568
rect 345164 7556 345170 7608
rect 371694 7556 371700 7608
rect 371752 7596 371758 7608
rect 436738 7596 436744 7608
rect 371752 7568 436744 7596
rect 371752 7556 371758 7568
rect 436738 7556 436744 7568
rect 436796 7556 436802 7608
rect 77386 7488 77392 7540
rect 77444 7528 77450 7540
rect 234706 7528 234712 7540
rect 77444 7500 234712 7528
rect 77444 7488 77450 7500
rect 234706 7488 234712 7500
rect 234764 7488 234770 7540
rect 101030 7420 101036 7472
rect 101088 7460 101094 7472
rect 251266 7460 251272 7472
rect 101088 7432 251272 7460
rect 101088 7420 101094 7432
rect 251266 7420 251272 7432
rect 251324 7420 251330 7472
rect 128170 7352 128176 7404
rect 128228 7392 128234 7404
rect 270494 7392 270500 7404
rect 128228 7364 270500 7392
rect 128228 7352 128234 7364
rect 270494 7352 270500 7364
rect 270552 7352 270558 7404
rect 158898 7284 158904 7336
rect 158956 7324 158962 7336
rect 291194 7324 291200 7336
rect 158956 7296 291200 7324
rect 158956 7284 158962 7296
rect 291194 7284 291200 7296
rect 291252 7284 291258 7336
rect 163682 7216 163688 7268
rect 163740 7256 163746 7268
rect 294046 7256 294052 7268
rect 163740 7228 294052 7256
rect 163740 7216 163746 7228
rect 294046 7216 294052 7228
rect 294104 7216 294110 7268
rect 167178 7148 167184 7200
rect 167236 7188 167242 7200
rect 296806 7188 296812 7200
rect 167236 7160 296812 7188
rect 167236 7148 167242 7160
rect 296806 7148 296812 7160
rect 296864 7148 296870 7200
rect 170766 7080 170772 7132
rect 170824 7120 170830 7132
rect 299566 7120 299572 7132
rect 170824 7092 299572 7120
rect 170824 7080 170830 7092
rect 299566 7080 299572 7092
rect 299624 7080 299630 7132
rect 174262 7012 174268 7064
rect 174320 7052 174326 7064
rect 302234 7052 302240 7064
rect 174320 7024 302240 7052
rect 174320 7012 174326 7024
rect 302234 7012 302240 7024
rect 302292 7012 302298 7064
rect 162486 6808 162492 6860
rect 162544 6848 162550 6860
rect 293954 6848 293960 6860
rect 162544 6820 293960 6848
rect 162544 6808 162550 6820
rect 293954 6808 293960 6820
rect 294012 6808 294018 6860
rect 130562 6740 130568 6792
rect 130620 6780 130626 6792
rect 271966 6780 271972 6792
rect 130620 6752 271972 6780
rect 130620 6740 130626 6752
rect 271966 6740 271972 6752
rect 272024 6740 272030 6792
rect 374086 6740 374092 6792
rect 374144 6780 374150 6792
rect 438854 6780 438860 6792
rect 374144 6752 438860 6780
rect 374144 6740 374150 6752
rect 438854 6740 438860 6752
rect 438912 6740 438918 6792
rect 126974 6672 126980 6724
rect 127032 6712 127038 6724
rect 269206 6712 269212 6724
rect 127032 6684 269212 6712
rect 127032 6672 127038 6684
rect 269206 6672 269212 6684
rect 269264 6672 269270 6724
rect 370682 6672 370688 6724
rect 370740 6712 370746 6724
rect 436186 6712 436192 6724
rect 370740 6684 436192 6712
rect 370740 6672 370746 6684
rect 436186 6672 436192 6684
rect 436244 6672 436250 6724
rect 97442 6604 97448 6656
rect 97500 6644 97506 6656
rect 248506 6644 248512 6656
rect 97500 6616 248512 6644
rect 97500 6604 97506 6616
rect 248506 6604 248512 6616
rect 248564 6604 248570 6656
rect 367002 6604 367008 6656
rect 367060 6644 367066 6656
rect 434714 6644 434720 6656
rect 367060 6616 434720 6644
rect 367060 6604 367066 6616
rect 434714 6604 434720 6616
rect 434772 6604 434778 6656
rect 93946 6536 93952 6588
rect 94004 6576 94010 6588
rect 247126 6576 247132 6588
rect 94004 6548 247132 6576
rect 94004 6536 94010 6548
rect 247126 6536 247132 6548
rect 247184 6536 247190 6588
rect 339862 6536 339868 6588
rect 339920 6576 339926 6588
rect 410518 6576 410524 6588
rect 339920 6548 410524 6576
rect 339920 6536 339926 6548
rect 410518 6536 410524 6548
rect 410576 6536 410582 6588
rect 90450 6468 90456 6520
rect 90508 6508 90514 6520
rect 244274 6508 244280 6520
rect 90508 6480 244280 6508
rect 90508 6468 90514 6480
rect 244274 6468 244280 6480
rect 244332 6468 244338 6520
rect 292574 6468 292580 6520
rect 292632 6508 292638 6520
rect 382366 6508 382372 6520
rect 292632 6480 382372 6508
rect 292632 6468 292638 6480
rect 382366 6468 382372 6480
rect 382424 6468 382430 6520
rect 86862 6400 86868 6452
rect 86920 6440 86926 6452
rect 241606 6440 241612 6452
rect 86920 6412 241612 6440
rect 86920 6400 86926 6412
rect 241606 6400 241612 6412
rect 241664 6400 241670 6452
rect 288986 6400 288992 6452
rect 289044 6440 289050 6452
rect 380894 6440 380900 6452
rect 289044 6412 380900 6440
rect 289044 6400 289050 6412
rect 380894 6400 380900 6412
rect 380952 6400 380958 6452
rect 389450 6400 389456 6452
rect 389508 6440 389514 6452
rect 449158 6440 449164 6452
rect 389508 6412 449164 6440
rect 389508 6400 389514 6412
rect 449158 6400 449164 6412
rect 449216 6400 449222 6452
rect 83274 6332 83280 6384
rect 83332 6372 83338 6384
rect 238846 6372 238852 6384
rect 83332 6344 238852 6372
rect 83332 6332 83338 6344
rect 238846 6332 238852 6344
rect 238904 6332 238910 6384
rect 285398 6332 285404 6384
rect 285456 6372 285462 6384
rect 378134 6372 378140 6384
rect 285456 6344 378140 6372
rect 285456 6332 285462 6344
rect 378134 6332 378140 6344
rect 378192 6332 378198 6384
rect 382366 6332 382372 6384
rect 382424 6372 382430 6384
rect 443638 6372 443644 6384
rect 382424 6344 443644 6372
rect 382424 6332 382430 6344
rect 443638 6332 443644 6344
rect 443696 6332 443702 6384
rect 79686 6264 79692 6316
rect 79744 6304 79750 6316
rect 237374 6304 237380 6316
rect 79744 6276 237380 6304
rect 79744 6264 79750 6276
rect 237374 6264 237380 6276
rect 237432 6264 237438 6316
rect 281902 6264 281908 6316
rect 281960 6304 281966 6316
rect 375466 6304 375472 6316
rect 281960 6276 375472 6304
rect 281960 6264 281966 6276
rect 375466 6264 375472 6276
rect 375524 6264 375530 6316
rect 384758 6264 384764 6316
rect 384816 6304 384822 6316
rect 445846 6304 445852 6316
rect 384816 6276 445852 6304
rect 384816 6264 384822 6276
rect 445846 6264 445852 6276
rect 445904 6264 445910 6316
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 187786 6236 187792 6248
rect 8812 6208 187792 6236
rect 8812 6196 8818 6208
rect 187786 6196 187792 6208
rect 187844 6196 187850 6248
rect 190822 6196 190828 6248
rect 190880 6236 190886 6248
rect 313366 6236 313372 6248
rect 190880 6208 313372 6236
rect 190880 6196 190886 6208
rect 313366 6196 313372 6208
rect 313424 6196 313430 6248
rect 346946 6196 346952 6248
rect 347004 6236 347010 6248
rect 421006 6236 421012 6248
rect 347004 6208 421012 6236
rect 347004 6196 347010 6208
rect 421006 6196 421012 6208
rect 421064 6196 421070 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 184934 6168 184940 6180
rect 4120 6140 184940 6168
rect 4120 6128 4126 6140
rect 184934 6128 184940 6140
rect 184992 6128 184998 6180
rect 187326 6128 187332 6180
rect 187384 6168 187390 6180
rect 310606 6168 310612 6180
rect 187384 6140 310612 6168
rect 187384 6128 187390 6140
rect 310606 6128 310612 6140
rect 310664 6128 310670 6180
rect 311618 6128 311624 6180
rect 311676 6168 311682 6180
rect 393406 6168 393412 6180
rect 311676 6140 393412 6168
rect 311676 6128 311682 6140
rect 393406 6128 393412 6140
rect 393464 6128 393470 6180
rect 501782 6128 501788 6180
rect 501840 6168 501846 6180
rect 525150 6168 525156 6180
rect 501840 6140 525156 6168
rect 501840 6128 501846 6140
rect 525150 6128 525156 6140
rect 525208 6128 525214 6180
rect 166074 6060 166080 6112
rect 166132 6100 166138 6112
rect 296714 6100 296720 6112
rect 166132 6072 296720 6100
rect 166132 6060 166138 6072
rect 296714 6060 296720 6072
rect 296772 6060 296778 6112
rect 169570 5992 169576 6044
rect 169628 6032 169634 6044
rect 298186 6032 298192 6044
rect 169628 6004 298192 6032
rect 169628 5992 169634 6004
rect 298186 5992 298192 6004
rect 298244 5992 298250 6044
rect 173158 5924 173164 5976
rect 173216 5964 173222 5976
rect 300854 5964 300860 5976
rect 173216 5936 300860 5964
rect 173216 5924 173222 5936
rect 300854 5924 300860 5936
rect 300912 5924 300918 5976
rect 176654 5856 176660 5908
rect 176712 5896 176718 5908
rect 303614 5896 303620 5908
rect 176712 5868 303620 5896
rect 176712 5856 176718 5868
rect 303614 5856 303620 5868
rect 303672 5856 303678 5908
rect 180242 5788 180248 5840
rect 180300 5828 180306 5840
rect 306374 5828 306380 5840
rect 180300 5800 306380 5828
rect 180300 5788 180306 5800
rect 306374 5788 306380 5800
rect 306432 5788 306438 5840
rect 183738 5720 183744 5772
rect 183796 5760 183802 5772
rect 307846 5760 307852 5772
rect 183796 5732 307852 5760
rect 183796 5720 183802 5732
rect 307846 5720 307852 5732
rect 307904 5720 307910 5772
rect 194410 5652 194416 5704
rect 194468 5692 194474 5704
rect 316034 5692 316040 5704
rect 194468 5664 316040 5692
rect 194468 5652 194474 5664
rect 316034 5652 316040 5664
rect 316092 5652 316098 5704
rect 197906 5584 197912 5636
rect 197964 5624 197970 5636
rect 317506 5624 317512 5636
rect 197964 5596 317512 5624
rect 197964 5584 197970 5596
rect 317506 5584 317512 5596
rect 317564 5584 317570 5636
rect 47854 5448 47860 5500
rect 47912 5488 47918 5500
rect 215294 5488 215300 5500
rect 47912 5460 215300 5488
rect 47912 5448 47918 5460
rect 215294 5448 215300 5460
rect 215352 5448 215358 5500
rect 306742 5448 306748 5500
rect 306800 5488 306806 5500
rect 393314 5488 393320 5500
rect 306800 5460 393320 5488
rect 306800 5448 306806 5460
rect 393314 5448 393320 5460
rect 393372 5448 393378 5500
rect 33594 5380 33600 5432
rect 33652 5420 33658 5432
rect 205634 5420 205640 5432
rect 33652 5392 205640 5420
rect 33652 5380 33658 5392
rect 205634 5380 205640 5392
rect 205692 5380 205698 5432
rect 303154 5380 303160 5432
rect 303212 5420 303218 5432
rect 390554 5420 390560 5432
rect 303212 5392 390560 5420
rect 303212 5380 303218 5392
rect 390554 5380 390560 5392
rect 390612 5380 390618 5432
rect 30098 5312 30104 5364
rect 30156 5352 30162 5364
rect 202874 5352 202880 5364
rect 30156 5324 202880 5352
rect 30156 5312 30162 5324
rect 202874 5312 202880 5324
rect 202932 5312 202938 5364
rect 299658 5312 299664 5364
rect 299716 5352 299722 5364
rect 387794 5352 387800 5364
rect 299716 5324 387800 5352
rect 299716 5312 299722 5324
rect 387794 5312 387800 5324
rect 387852 5312 387858 5364
rect 26510 5244 26516 5296
rect 26568 5284 26574 5296
rect 200206 5284 200212 5296
rect 26568 5256 200212 5284
rect 26568 5244 26574 5256
rect 200206 5244 200212 5256
rect 200264 5244 200270 5296
rect 231394 5244 231400 5296
rect 231452 5284 231458 5296
rect 339494 5284 339500 5296
rect 231452 5256 339500 5284
rect 231452 5244 231458 5256
rect 339494 5244 339500 5256
rect 339552 5244 339558 5296
rect 342162 5244 342168 5296
rect 342220 5284 342226 5296
rect 416866 5284 416872 5296
rect 342220 5256 416872 5284
rect 342220 5244 342226 5256
rect 416866 5244 416872 5256
rect 416924 5244 416930 5296
rect 17034 5176 17040 5228
rect 17092 5216 17098 5228
rect 193306 5216 193312 5228
rect 17092 5188 193312 5216
rect 17092 5176 17098 5188
rect 193306 5176 193312 5188
rect 193364 5176 193370 5228
rect 215662 5176 215668 5228
rect 215720 5216 215726 5228
rect 329834 5216 329840 5228
rect 215720 5188 329840 5216
rect 215720 5176 215726 5188
rect 329834 5176 329840 5188
rect 329892 5176 329898 5228
rect 335078 5176 335084 5228
rect 335136 5216 335142 5228
rect 412634 5216 412640 5228
rect 335136 5188 412640 5216
rect 335136 5176 335142 5188
rect 412634 5176 412640 5188
rect 412692 5176 412698 5228
rect 21818 5108 21824 5160
rect 21876 5148 21882 5160
rect 197354 5148 197360 5160
rect 21876 5120 197360 5148
rect 21876 5108 21882 5120
rect 197354 5108 197360 5120
rect 197412 5108 197418 5160
rect 212534 5108 212540 5160
rect 212592 5148 212598 5160
rect 327074 5148 327080 5160
rect 212592 5120 327080 5148
rect 212592 5108 212598 5120
rect 327074 5108 327080 5120
rect 327132 5108 327138 5160
rect 331582 5108 331588 5160
rect 331640 5148 331646 5160
rect 409874 5148 409880 5160
rect 331640 5120 409880 5148
rect 331640 5108 331646 5120
rect 409874 5108 409880 5120
rect 409932 5108 409938 5160
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 190546 5080 190552 5092
rect 12400 5052 190552 5080
rect 12400 5040 12406 5052
rect 190546 5040 190552 5052
rect 190604 5040 190610 5092
rect 201494 5040 201500 5092
rect 201552 5080 201558 5092
rect 320174 5080 320180 5092
rect 201552 5052 320180 5080
rect 201552 5040 201558 5052
rect 320174 5040 320180 5052
rect 320232 5040 320238 5092
rect 320910 5040 320916 5092
rect 320968 5080 320974 5092
rect 402974 5080 402980 5092
rect 320968 5052 402980 5080
rect 320968 5040 320974 5052
rect 402974 5040 402980 5052
rect 403032 5040 403038 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 187694 5012 187700 5024
rect 7708 4984 187700 5012
rect 7708 4972 7714 4984
rect 187694 4972 187700 4984
rect 187752 4972 187758 5024
rect 205082 4972 205088 5024
rect 205140 5012 205146 5024
rect 322934 5012 322940 5024
rect 205140 4984 322940 5012
rect 205140 4972 205146 4984
rect 322934 4972 322940 4984
rect 322992 4972 322998 5024
rect 324406 4972 324412 5024
rect 324464 5012 324470 5024
rect 404446 5012 404452 5024
rect 324464 4984 404452 5012
rect 324464 4972 324470 4984
rect 404446 4972 404452 4984
rect 404504 4972 404510 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 183554 4944 183560 4956
rect 2924 4916 183560 4944
rect 2924 4904 2930 4916
rect 183554 4904 183560 4916
rect 183612 4904 183618 4956
rect 202690 4904 202696 4956
rect 202748 4944 202754 4956
rect 321554 4944 321560 4956
rect 202748 4916 321560 4944
rect 202748 4904 202754 4916
rect 321554 4904 321560 4916
rect 321612 4904 321618 4956
rect 327994 4904 328000 4956
rect 328052 4944 328058 4956
rect 407206 4944 407212 4956
rect 328052 4916 407212 4944
rect 328052 4904 328058 4916
rect 407206 4904 407212 4916
rect 407264 4904 407270 4956
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 182174 4876 182180 4888
rect 624 4848 182180 4876
rect 624 4836 630 4848
rect 182174 4836 182180 4848
rect 182232 4836 182238 4888
rect 192018 4836 192024 4888
rect 192076 4876 192082 4888
rect 313274 4876 313280 4888
rect 192076 4848 313280 4876
rect 192076 4836 192082 4848
rect 313274 4836 313280 4848
rect 313332 4836 313338 4888
rect 313826 4836 313832 4888
rect 313884 4876 313890 4888
rect 397454 4876 397460 4888
rect 313884 4848 397460 4876
rect 313884 4836 313890 4848
rect 397454 4836 397460 4848
rect 397512 4836 397518 4888
rect 459186 4836 459192 4888
rect 459244 4876 459250 4888
rect 496906 4876 496912 4888
rect 459244 4848 496912 4876
rect 459244 4836 459250 4848
rect 496906 4836 496912 4848
rect 496964 4836 496970 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 183646 4808 183652 4820
rect 1728 4780 183652 4808
rect 1728 4768 1734 4780
rect 183646 4768 183652 4780
rect 183704 4768 183710 4820
rect 184934 4768 184940 4820
rect 184992 4808 184998 4820
rect 309134 4808 309140 4820
rect 184992 4780 309140 4808
rect 184992 4768 184998 4780
rect 309134 4768 309140 4780
rect 309192 4768 309198 4820
rect 310238 4768 310244 4820
rect 310296 4808 310302 4820
rect 394786 4808 394792 4820
rect 310296 4780 394792 4808
rect 310296 4768 310302 4780
rect 394786 4768 394792 4780
rect 394844 4768 394850 4820
rect 420178 4768 420184 4820
rect 420236 4808 420242 4820
rect 470594 4808 470600 4820
rect 420236 4780 470600 4808
rect 420236 4768 420242 4780
rect 470594 4768 470600 4780
rect 470652 4768 470658 4820
rect 51350 4700 51356 4752
rect 51408 4740 51414 4752
rect 218054 4740 218060 4752
rect 51408 4712 218060 4740
rect 51408 4700 51414 4712
rect 218054 4700 218060 4712
rect 218112 4700 218118 4752
rect 317322 4700 317328 4752
rect 317380 4740 317386 4752
rect 400214 4740 400220 4752
rect 317380 4712 400220 4740
rect 317380 4700 317386 4712
rect 400214 4700 400220 4712
rect 400272 4700 400278 4752
rect 54938 4632 54944 4684
rect 54996 4672 55002 4684
rect 219526 4672 219532 4684
rect 54996 4644 219532 4672
rect 54996 4632 55002 4644
rect 219526 4632 219532 4644
rect 219584 4632 219590 4684
rect 338666 4632 338672 4684
rect 338724 4672 338730 4684
rect 414106 4672 414112 4684
rect 338724 4644 414112 4672
rect 338724 4632 338730 4644
rect 414106 4632 414112 4644
rect 414164 4632 414170 4684
rect 62022 4564 62028 4616
rect 62080 4604 62086 4616
rect 224954 4604 224960 4616
rect 62080 4576 224960 4604
rect 62080 4564 62086 4576
rect 224954 4564 224960 4576
rect 225012 4564 225018 4616
rect 345750 4564 345756 4616
rect 345808 4604 345814 4616
rect 419534 4604 419540 4616
rect 345808 4576 419540 4604
rect 345808 4564 345814 4576
rect 419534 4564 419540 4576
rect 419592 4564 419598 4616
rect 58434 4496 58440 4548
rect 58492 4536 58498 4548
rect 222194 4536 222200 4548
rect 58492 4508 222200 4536
rect 58492 4496 58498 4508
rect 222194 4496 222200 4508
rect 222252 4496 222258 4548
rect 349246 4496 349252 4548
rect 349304 4536 349310 4548
rect 422294 4536 422300 4548
rect 349304 4508 422300 4536
rect 349304 4496 349310 4508
rect 422294 4496 422300 4508
rect 422352 4496 422358 4548
rect 65518 4428 65524 4480
rect 65576 4468 65582 4480
rect 227714 4468 227720 4480
rect 65576 4440 227720 4468
rect 65576 4428 65582 4440
rect 227714 4428 227720 4440
rect 227772 4428 227778 4480
rect 352834 4428 352840 4480
rect 352892 4468 352898 4480
rect 423766 4468 423772 4480
rect 352892 4440 423772 4468
rect 352892 4428 352898 4440
rect 423766 4428 423772 4440
rect 423824 4428 423830 4480
rect 72602 4360 72608 4412
rect 72660 4400 72666 4412
rect 231946 4400 231952 4412
rect 72660 4372 231952 4400
rect 72660 4360 72666 4372
rect 231946 4360 231952 4372
rect 232004 4360 232010 4412
rect 356330 4360 356336 4412
rect 356388 4400 356394 4412
rect 426526 4400 426532 4412
rect 356388 4372 426532 4400
rect 356388 4360 356394 4372
rect 426526 4360 426532 4372
rect 426584 4360 426590 4412
rect 69106 4292 69112 4344
rect 69164 4332 69170 4344
rect 229186 4332 229192 4344
rect 69164 4304 229192 4332
rect 69164 4292 69170 4304
rect 229186 4292 229192 4304
rect 229244 4292 229250 4344
rect 359918 4292 359924 4344
rect 359976 4332 359982 4344
rect 429194 4332 429200 4344
rect 359976 4304 429200 4332
rect 359976 4292 359982 4304
rect 429194 4292 429200 4304
rect 429252 4292 429258 4344
rect 76190 4224 76196 4276
rect 76248 4264 76254 4276
rect 234614 4264 234620 4276
rect 76248 4236 234620 4264
rect 76248 4224 76254 4236
rect 234614 4224 234620 4236
rect 234672 4224 234678 4276
rect 363506 4224 363512 4276
rect 363564 4264 363570 4276
rect 431954 4264 431960 4276
rect 363564 4236 431960 4264
rect 363564 4224 363570 4236
rect 431954 4224 431960 4236
rect 432012 4224 432018 4276
rect 486344 4168 486556 4196
rect 67910 4088 67916 4140
rect 67968 4128 67974 4140
rect 214650 4128 214656 4140
rect 67968 4100 214656 4128
rect 67968 4088 67974 4100
rect 214650 4088 214656 4100
rect 214708 4088 214714 4140
rect 226334 4088 226340 4140
rect 226392 4128 226398 4140
rect 256050 4128 256056 4140
rect 226392 4100 256056 4128
rect 226392 4088 226398 4100
rect 256050 4088 256056 4100
rect 256108 4088 256114 4140
rect 258166 4088 258172 4140
rect 258224 4128 258230 4140
rect 258718 4128 258724 4140
rect 258224 4100 258724 4128
rect 258224 4088 258230 4100
rect 258718 4088 258724 4100
rect 258776 4088 258782 4140
rect 259454 4088 259460 4140
rect 259512 4128 259518 4140
rect 305454 4128 305460 4140
rect 259512 4100 305460 4128
rect 259512 4088 259518 4100
rect 305454 4088 305460 4100
rect 305512 4088 305518 4140
rect 319714 4088 319720 4140
rect 319772 4128 319778 4140
rect 399478 4128 399484 4140
rect 319772 4100 399484 4128
rect 319772 4088 319778 4100
rect 399478 4088 399484 4100
rect 399536 4088 399542 4140
rect 402514 4088 402520 4140
rect 402572 4128 402578 4140
rect 403526 4128 403532 4140
rect 402572 4100 403532 4128
rect 402572 4088 402578 4100
rect 403526 4088 403532 4100
rect 403584 4088 403590 4140
rect 416593 4131 416651 4137
rect 416593 4097 416605 4131
rect 416639 4128 416651 4131
rect 463694 4128 463700 4140
rect 416639 4100 463700 4128
rect 416639 4097 416651 4100
rect 416593 4091 416651 4097
rect 463694 4088 463700 4100
rect 463752 4088 463758 4140
rect 469214 4128 469220 4140
rect 463896 4100 469220 4128
rect 28813 4063 28871 4069
rect 28813 4029 28825 4063
rect 28859 4060 28871 4063
rect 35158 4060 35164 4072
rect 28859 4032 35164 4060
rect 28859 4029 28871 4032
rect 28813 4023 28871 4029
rect 35158 4020 35164 4032
rect 35216 4020 35222 4072
rect 38378 4020 38384 4072
rect 38436 4060 38442 4072
rect 47578 4060 47584 4072
rect 38436 4032 47584 4060
rect 38436 4020 38442 4032
rect 47578 4020 47584 4032
rect 47636 4020 47642 4072
rect 50065 4063 50123 4069
rect 50065 4029 50077 4063
rect 50111 4060 50123 4063
rect 57238 4060 57244 4072
rect 50111 4032 57244 4060
rect 50111 4029 50123 4032
rect 50065 4023 50123 4029
rect 57238 4020 57244 4032
rect 57296 4020 57302 4072
rect 60826 4020 60832 4072
rect 60884 4060 60890 4072
rect 204901 4063 204959 4069
rect 204901 4060 204913 4063
rect 60884 4032 204913 4060
rect 60884 4020 60890 4032
rect 204901 4029 204913 4032
rect 204947 4029 204959 4063
rect 204901 4023 204959 4029
rect 221550 4020 221556 4072
rect 221608 4060 221614 4072
rect 253382 4060 253388 4072
rect 221608 4032 253388 4060
rect 221608 4020 221614 4032
rect 253382 4020 253388 4032
rect 253440 4020 253446 4072
rect 257062 4020 257068 4072
rect 257120 4060 257126 4072
rect 271138 4060 271144 4072
rect 257120 4032 271144 4060
rect 257120 4020 257126 4032
rect 271138 4020 271144 4032
rect 271196 4020 271202 4072
rect 298462 4020 298468 4072
rect 298520 4060 298526 4072
rect 378781 4063 378839 4069
rect 378781 4060 378793 4063
rect 298520 4032 378793 4060
rect 298520 4020 298526 4032
rect 378781 4029 378793 4032
rect 378827 4029 378839 4063
rect 378781 4023 378839 4029
rect 403618 4020 403624 4072
rect 403676 4060 403682 4072
rect 459738 4060 459744 4072
rect 403676 4032 459744 4060
rect 403676 4020 403682 4032
rect 459738 4020 459744 4032
rect 459796 4020 459802 4072
rect 462593 4063 462651 4069
rect 462593 4029 462605 4063
rect 462639 4060 462651 4063
rect 463896 4060 463924 4100
rect 469214 4088 469220 4100
rect 469272 4088 469278 4140
rect 469858 4088 469864 4140
rect 469916 4128 469922 4140
rect 471238 4128 471244 4140
rect 469916 4100 471244 4128
rect 469916 4088 469922 4100
rect 471238 4088 471244 4100
rect 471296 4088 471302 4140
rect 485041 4131 485099 4137
rect 485041 4128 485053 4131
rect 471992 4100 485053 4128
rect 462639 4032 463924 4060
rect 462639 4029 462651 4032
rect 462593 4023 462651 4029
rect 468662 4020 468668 4072
rect 468720 4060 468726 4072
rect 471992 4060 472020 4100
rect 485041 4097 485053 4100
rect 485087 4097 485099 4131
rect 485041 4091 485099 4097
rect 468720 4032 472020 4060
rect 468720 4020 468726 4032
rect 475746 4020 475752 4072
rect 475804 4060 475810 4072
rect 486344 4060 486372 4168
rect 486528 4128 486556 4168
rect 486528 4100 489914 4128
rect 475804 4032 486372 4060
rect 489886 4060 489914 4100
rect 505370 4088 505376 4140
rect 505428 4128 505434 4140
rect 511166 4128 511172 4140
rect 505428 4100 511172 4128
rect 505428 4088 505434 4100
rect 511166 4088 511172 4100
rect 511224 4088 511230 4140
rect 500218 4060 500224 4072
rect 489886 4032 500224 4060
rect 475804 4020 475810 4032
rect 500218 4020 500224 4032
rect 500276 4020 500282 4072
rect 524230 4020 524236 4072
rect 524288 4060 524294 4072
rect 529198 4060 529204 4072
rect 524288 4032 529204 4060
rect 524288 4020 524294 4032
rect 529198 4020 529204 4032
rect 529256 4020 529262 4072
rect 14734 3952 14740 4004
rect 14792 3992 14798 4004
rect 18598 3992 18604 4004
rect 14792 3964 18604 3992
rect 14792 3952 14798 3964
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 34790 3952 34796 4004
rect 34848 3992 34854 4004
rect 51810 3992 51816 4004
rect 34848 3964 51816 3992
rect 34848 3952 34854 3964
rect 51810 3952 51816 3964
rect 51868 3952 51874 4004
rect 53742 3952 53748 4004
rect 53800 3992 53806 4004
rect 210418 3992 210424 4004
rect 53800 3964 210424 3992
rect 53800 3952 53806 3964
rect 210418 3952 210424 3964
rect 210476 3952 210482 4004
rect 219250 3952 219256 4004
rect 219308 3992 219314 4004
rect 251818 3992 251824 4004
rect 219308 3964 251824 3992
rect 219308 3952 219314 3964
rect 251818 3952 251824 3964
rect 251876 3952 251882 4004
rect 254670 3952 254676 4004
rect 254728 3992 254734 4004
rect 273898 3992 273904 4004
rect 254728 3964 273904 3992
rect 254728 3952 254734 3964
rect 273898 3952 273904 3964
rect 273956 3952 273962 4004
rect 276014 3952 276020 4004
rect 276072 3992 276078 4004
rect 291838 3992 291844 4004
rect 276072 3964 291844 3992
rect 276072 3952 276078 3964
rect 291838 3952 291844 3964
rect 291896 3952 291902 4004
rect 293678 3952 293684 4004
rect 293736 3992 293742 4004
rect 298738 3992 298744 4004
rect 293736 3964 298744 3992
rect 293736 3952 293742 3964
rect 298738 3952 298744 3964
rect 298796 3952 298802 4004
rect 305546 3952 305552 4004
rect 305604 3992 305610 4004
rect 391198 3992 391204 4004
rect 305604 3964 391204 3992
rect 305604 3952 305610 3964
rect 391198 3952 391204 3964
rect 391256 3952 391262 4004
rect 393038 3952 393044 4004
rect 393096 3992 393102 4004
rect 396810 3992 396816 4004
rect 393096 3964 396816 3992
rect 393096 3952 393102 3964
rect 396810 3952 396816 3964
rect 396868 3952 396874 4004
rect 397730 3952 397736 4004
rect 397788 3992 397794 4004
rect 455414 3992 455420 4004
rect 397788 3964 455420 3992
rect 397788 3952 397794 3964
rect 455414 3952 455420 3964
rect 455472 3952 455478 4004
rect 460382 3952 460388 4004
rect 460440 3992 460446 4004
rect 486326 3992 486332 4004
rect 460440 3964 486332 3992
rect 460440 3952 460446 3964
rect 486326 3952 486332 3964
rect 486384 3952 486390 4004
rect 25314 3884 25320 3936
rect 25372 3924 25378 3936
rect 29638 3924 29644 3936
rect 25372 3896 29644 3924
rect 25372 3884 25378 3896
rect 29638 3884 29644 3896
rect 29696 3884 29702 3936
rect 31294 3884 31300 3936
rect 31352 3924 31358 3936
rect 39298 3924 39304 3936
rect 31352 3896 39304 3924
rect 31352 3884 31358 3896
rect 39298 3884 39304 3896
rect 39356 3884 39362 3936
rect 43070 3884 43076 3936
rect 43128 3924 43134 3936
rect 204809 3927 204867 3933
rect 204809 3924 204821 3927
rect 43128 3896 204821 3924
rect 43128 3884 43134 3896
rect 204809 3893 204821 3896
rect 204855 3893 204867 3927
rect 204809 3887 204867 3893
rect 204901 3927 204959 3933
rect 204901 3893 204913 3927
rect 204947 3924 204959 3927
rect 211798 3924 211804 3936
rect 204947 3896 211804 3924
rect 204947 3893 204959 3896
rect 204901 3887 204959 3893
rect 211798 3884 211804 3896
rect 211856 3884 211862 3936
rect 225138 3884 225144 3936
rect 225196 3924 225202 3936
rect 264238 3924 264244 3936
rect 225196 3896 264244 3924
rect 225196 3884 225202 3896
rect 264238 3884 264244 3896
rect 264296 3884 264302 3936
rect 266538 3884 266544 3936
rect 266596 3924 266602 3936
rect 268378 3924 268384 3936
rect 266596 3896 268384 3924
rect 266596 3884 266602 3896
rect 268378 3884 268384 3896
rect 268436 3884 268442 3936
rect 272426 3884 272432 3936
rect 272484 3924 272490 3936
rect 279421 3927 279479 3933
rect 279421 3924 279433 3927
rect 272484 3896 279433 3924
rect 272484 3884 272490 3896
rect 279421 3893 279433 3896
rect 279467 3893 279479 3927
rect 279421 3887 279479 3893
rect 279510 3884 279516 3936
rect 279568 3924 279574 3936
rect 289078 3924 289084 3936
rect 279568 3896 289084 3924
rect 279568 3884 279574 3896
rect 289078 3884 289084 3896
rect 289136 3884 289142 3936
rect 297177 3927 297235 3933
rect 297177 3893 297189 3927
rect 297223 3924 297235 3927
rect 382274 3924 382280 3936
rect 297223 3896 382280 3924
rect 297223 3893 297235 3896
rect 297177 3887 297235 3893
rect 382274 3884 382280 3896
rect 382332 3884 382338 3936
rect 388073 3927 388131 3933
rect 388073 3893 388085 3927
rect 388119 3924 388131 3927
rect 392578 3924 392584 3936
rect 388119 3896 392584 3924
rect 388119 3893 388131 3896
rect 388073 3887 388131 3893
rect 392578 3884 392584 3896
rect 392636 3884 392642 3936
rect 404081 3927 404139 3933
rect 404081 3893 404093 3927
rect 404127 3924 404139 3927
rect 454034 3924 454040 3936
rect 404127 3896 454040 3924
rect 404127 3893 404139 3896
rect 404081 3887 404139 3893
rect 454034 3884 454040 3896
rect 454092 3884 454098 3936
rect 454494 3884 454500 3936
rect 454552 3924 454558 3936
rect 480898 3924 480904 3936
rect 454552 3896 480904 3924
rect 454552 3884 454558 3896
rect 480898 3884 480904 3896
rect 480956 3884 480962 3936
rect 485041 3927 485099 3933
rect 485041 3893 485053 3927
rect 485087 3924 485099 3927
rect 492030 3924 492036 3936
rect 485087 3896 492036 3924
rect 485087 3893 485099 3896
rect 485041 3887 485099 3893
rect 492030 3884 492036 3896
rect 492088 3884 492094 3936
rect 504174 3884 504180 3936
rect 504232 3924 504238 3936
rect 522298 3924 522304 3936
rect 504232 3896 522304 3924
rect 504232 3884 504238 3896
rect 522298 3884 522304 3896
rect 522356 3884 522362 3936
rect 24210 3816 24216 3868
rect 24268 3856 24274 3868
rect 28813 3859 28871 3865
rect 28813 3856 28825 3859
rect 24268 3828 28825 3856
rect 24268 3816 24274 3828
rect 28813 3825 28825 3828
rect 28859 3825 28871 3859
rect 28813 3819 28871 3825
rect 28902 3816 28908 3868
rect 28960 3856 28966 3868
rect 28960 3828 35894 3856
rect 28960 3816 28966 3828
rect 27706 3748 27712 3800
rect 27764 3788 27770 3800
rect 32398 3788 32404 3800
rect 27764 3760 32404 3788
rect 27764 3748 27770 3760
rect 32398 3748 32404 3760
rect 32456 3748 32462 3800
rect 35866 3788 35894 3828
rect 35986 3816 35992 3868
rect 36044 3856 36050 3868
rect 207014 3856 207020 3868
rect 36044 3828 207020 3856
rect 36044 3816 36050 3828
rect 207014 3816 207020 3828
rect 207072 3816 207078 3868
rect 234614 3816 234620 3868
rect 234672 3856 234678 3868
rect 240778 3856 240784 3868
rect 234672 3828 240784 3856
rect 234672 3816 234678 3828
rect 240778 3816 240784 3828
rect 240836 3816 240842 3868
rect 241609 3859 241667 3865
rect 241609 3825 241621 3859
rect 241655 3856 241667 3859
rect 274082 3856 274088 3868
rect 241655 3828 274088 3856
rect 241655 3825 241667 3828
rect 241609 3819 241667 3825
rect 274082 3816 274088 3828
rect 274140 3816 274146 3868
rect 284294 3816 284300 3868
rect 284352 3856 284358 3868
rect 376754 3856 376760 3868
rect 284352 3828 376760 3856
rect 284352 3816 284358 3828
rect 376754 3816 376760 3828
rect 376812 3816 376818 3868
rect 378781 3859 378839 3865
rect 378781 3825 378793 3859
rect 378827 3856 378839 3859
rect 384298 3856 384304 3868
rect 378827 3828 384304 3856
rect 378827 3825 378839 3828
rect 378781 3819 378839 3825
rect 384298 3816 384304 3828
rect 384356 3816 384362 3868
rect 390646 3816 390652 3868
rect 390704 3856 390710 3868
rect 449986 3856 449992 3868
rect 390704 3828 449992 3856
rect 390704 3816 390710 3828
rect 449986 3816 449992 3828
rect 450044 3816 450050 3868
rect 461578 3816 461584 3868
rect 461636 3856 461642 3868
rect 491938 3856 491944 3868
rect 461636 3828 491944 3856
rect 461636 3816 461642 3828
rect 491938 3816 491944 3828
rect 491996 3816 492002 3868
rect 497090 3816 497096 3868
rect 497148 3856 497154 3868
rect 519446 3856 519452 3868
rect 497148 3828 519452 3856
rect 497148 3816 497154 3828
rect 519446 3816 519452 3828
rect 519504 3816 519510 3868
rect 531314 3816 531320 3868
rect 531372 3856 531378 3868
rect 546678 3856 546684 3868
rect 531372 3828 546684 3856
rect 531372 3816 531378 3828
rect 546678 3816 546684 3828
rect 546736 3816 546742 3868
rect 204809 3791 204867 3797
rect 35866 3760 200114 3788
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 195974 3720 195980 3732
rect 20680 3692 195980 3720
rect 20680 3680 20686 3692
rect 195974 3680 195980 3692
rect 196032 3680 196038 3732
rect 200086 3720 200114 3760
rect 204809 3757 204821 3791
rect 204855 3788 204867 3791
rect 211154 3788 211160 3800
rect 204855 3760 211160 3788
rect 204855 3757 204867 3760
rect 204809 3751 204867 3757
rect 211154 3748 211160 3760
rect 211212 3748 211218 3800
rect 214466 3748 214472 3800
rect 214524 3788 214530 3800
rect 258077 3791 258135 3797
rect 258077 3788 258089 3791
rect 214524 3760 258089 3788
rect 214524 3748 214530 3760
rect 258077 3757 258089 3760
rect 258123 3757 258135 3791
rect 262858 3788 262864 3800
rect 258077 3751 258135 3757
rect 258184 3760 262864 3788
rect 201586 3720 201592 3732
rect 200086 3692 201592 3720
rect 201586 3680 201592 3692
rect 201644 3680 201650 3732
rect 210970 3680 210976 3732
rect 211028 3720 211034 3732
rect 258184 3720 258212 3760
rect 262858 3748 262864 3760
rect 262916 3748 262922 3800
rect 270034 3748 270040 3800
rect 270092 3788 270098 3800
rect 270092 3760 271920 3788
rect 270092 3748 270098 3760
rect 211028 3692 258212 3720
rect 211028 3680 211034 3692
rect 263042 3680 263048 3732
rect 263100 3720 263106 3732
rect 263100 3692 267228 3720
rect 263100 3680 263106 3692
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 196066 3652 196072 3664
rect 19484 3624 196072 3652
rect 19484 3612 19490 3624
rect 196066 3612 196072 3624
rect 196124 3612 196130 3664
rect 207382 3612 207388 3664
rect 207440 3652 207446 3664
rect 258166 3652 258172 3664
rect 207440 3624 258172 3652
rect 207440 3612 207446 3624
rect 258166 3612 258172 3624
rect 258224 3612 258230 3664
rect 258258 3612 258264 3664
rect 258316 3652 258322 3664
rect 259362 3652 259368 3664
rect 258316 3624 259368 3652
rect 258316 3612 258322 3624
rect 259362 3612 259368 3624
rect 259420 3612 259426 3664
rect 261754 3612 261760 3664
rect 261812 3652 261818 3664
rect 262950 3652 262956 3664
rect 261812 3624 262956 3652
rect 261812 3612 261818 3624
rect 262950 3612 262956 3624
rect 263008 3612 263014 3664
rect 264146 3612 264152 3664
rect 264204 3652 264210 3664
rect 264882 3652 264888 3664
rect 264204 3624 264888 3652
rect 264204 3612 264210 3624
rect 264882 3612 264888 3624
rect 264940 3612 264946 3664
rect 265342 3612 265348 3664
rect 265400 3652 265406 3664
rect 267090 3652 267096 3664
rect 265400 3624 267096 3652
rect 265400 3612 265406 3624
rect 267090 3612 267096 3624
rect 267148 3612 267154 3664
rect 267200 3652 267228 3692
rect 267734 3680 267740 3732
rect 267792 3720 267798 3732
rect 269758 3720 269764 3732
rect 267792 3692 269764 3720
rect 267792 3680 267798 3692
rect 269758 3680 269764 3692
rect 269816 3680 269822 3732
rect 271230 3680 271236 3732
rect 271288 3720 271294 3732
rect 271782 3720 271788 3732
rect 271288 3692 271788 3720
rect 271288 3680 271294 3692
rect 271782 3680 271788 3692
rect 271840 3680 271846 3732
rect 271892 3720 271920 3760
rect 277118 3748 277124 3800
rect 277176 3788 277182 3800
rect 371878 3788 371884 3800
rect 277176 3760 371884 3788
rect 277176 3748 277182 3760
rect 371878 3748 371884 3760
rect 371936 3748 371942 3800
rect 378870 3748 378876 3800
rect 378928 3788 378934 3800
rect 380158 3788 380164 3800
rect 378928 3760 380164 3788
rect 378928 3748 378934 3760
rect 380158 3748 380164 3760
rect 380216 3748 380222 3800
rect 383562 3748 383568 3800
rect 383620 3788 383626 3800
rect 431957 3791 432015 3797
rect 431957 3788 431969 3791
rect 383620 3760 431969 3788
rect 383620 3748 383626 3760
rect 431957 3757 431969 3760
rect 432003 3757 432015 3791
rect 431957 3751 432015 3757
rect 432046 3748 432052 3800
rect 432104 3788 432110 3800
rect 432104 3760 440372 3788
rect 432104 3748 432110 3760
rect 367094 3720 367100 3732
rect 271892 3692 367100 3720
rect 367094 3680 367100 3692
rect 367152 3680 367158 3732
rect 369394 3680 369400 3732
rect 369452 3720 369458 3732
rect 369452 3692 370728 3720
rect 369452 3680 369458 3692
rect 355137 3655 355195 3661
rect 355137 3652 355149 3655
rect 267200 3624 355149 3652
rect 355137 3621 355149 3624
rect 355183 3621 355195 3655
rect 355137 3615 355195 3621
rect 355226 3612 355232 3664
rect 355284 3652 355290 3664
rect 363693 3655 363751 3661
rect 363693 3652 363705 3655
rect 355284 3624 363705 3652
rect 355284 3612 355290 3624
rect 363693 3621 363705 3624
rect 363739 3621 363751 3655
rect 363693 3615 363751 3621
rect 365806 3612 365812 3664
rect 365864 3652 365870 3664
rect 367738 3652 367744 3664
rect 365864 3624 367744 3652
rect 365864 3612 365870 3624
rect 367738 3612 367744 3624
rect 367796 3612 367802 3664
rect 368198 3612 368204 3664
rect 368256 3652 368262 3664
rect 370590 3652 370596 3664
rect 368256 3624 370596 3652
rect 368256 3612 368262 3624
rect 370590 3612 370596 3624
rect 370648 3612 370654 3664
rect 370700 3652 370728 3692
rect 372890 3680 372896 3732
rect 372948 3720 372954 3732
rect 373902 3720 373908 3732
rect 372948 3692 373908 3720
rect 372948 3680 372954 3692
rect 373902 3680 373908 3692
rect 373960 3680 373966 3732
rect 379974 3680 379980 3732
rect 380032 3720 380038 3732
rect 380802 3720 380808 3732
rect 380032 3692 380808 3720
rect 380032 3680 380038 3692
rect 380802 3680 380808 3692
rect 380860 3680 380866 3732
rect 381170 3680 381176 3732
rect 381228 3720 381234 3732
rect 382182 3720 382188 3732
rect 381228 3692 382188 3720
rect 381228 3680 381234 3692
rect 382182 3680 382188 3692
rect 382240 3680 382246 3732
rect 382277 3723 382335 3729
rect 382277 3689 382289 3723
rect 382323 3720 382335 3723
rect 436097 3723 436155 3729
rect 382323 3692 433104 3720
rect 382323 3689 382335 3692
rect 382277 3683 382335 3689
rect 370700 3624 433012 3652
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 11204 3556 190454 3584
rect 11204 3544 11210 3556
rect 190426 3528 190454 3556
rect 203886 3544 203892 3596
rect 203944 3584 203950 3596
rect 203944 3556 248414 3584
rect 203944 3544 203950 3556
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14458 3516 14464 3528
rect 13596 3488 14464 3516
rect 13596 3476 13602 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 181349 3519 181407 3525
rect 181349 3516 181361 3519
rect 14568 3488 181361 3516
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 5316 3420 9904 3448
rect 5316 3408 5322 3420
rect 6454 3272 6460 3324
rect 6512 3312 6518 3324
rect 7558 3312 7564 3324
rect 6512 3284 7564 3312
rect 6512 3272 6518 3284
rect 7558 3272 7564 3284
rect 7616 3272 7622 3324
rect 9876 3312 9904 3420
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 14568 3380 14596 3488
rect 181349 3485 181361 3488
rect 181395 3485 181407 3519
rect 181349 3479 181407 3485
rect 181438 3476 181444 3528
rect 181496 3516 181502 3528
rect 182082 3516 182088 3528
rect 181496 3488 182088 3516
rect 181496 3476 181502 3488
rect 182082 3476 182088 3488
rect 182140 3476 182146 3528
rect 182542 3476 182548 3528
rect 182600 3516 182606 3528
rect 183462 3516 183468 3528
rect 182600 3488 183468 3516
rect 182600 3476 182606 3488
rect 183462 3476 183468 3488
rect 183520 3476 183526 3528
rect 188522 3476 188528 3528
rect 188580 3516 188586 3528
rect 188982 3516 188988 3528
rect 188580 3488 188988 3516
rect 188580 3476 188586 3488
rect 188982 3476 188988 3488
rect 189040 3476 189046 3528
rect 190426 3488 190460 3528
rect 190454 3476 190460 3488
rect 190512 3476 190518 3528
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 194502 3516 194508 3528
rect 193272 3488 194508 3516
rect 193272 3476 193278 3488
rect 194502 3476 194508 3488
rect 194560 3476 194566 3528
rect 196802 3476 196808 3528
rect 196860 3516 196866 3528
rect 197262 3516 197268 3528
rect 196860 3488 197268 3516
rect 196860 3476 196866 3488
rect 197262 3476 197268 3488
rect 197320 3476 197326 3528
rect 208578 3476 208584 3528
rect 208636 3516 208642 3528
rect 209682 3516 209688 3528
rect 208636 3488 209688 3516
rect 208636 3476 208642 3488
rect 209682 3476 209688 3488
rect 209740 3476 209746 3528
rect 218054 3476 218060 3528
rect 218112 3516 218118 3528
rect 246298 3516 246304 3528
rect 218112 3488 246304 3516
rect 218112 3476 218118 3488
rect 246298 3476 246304 3488
rect 246356 3476 246362 3528
rect 248386 3516 248414 3556
rect 248782 3544 248788 3596
rect 248840 3584 248846 3596
rect 248840 3556 251220 3584
rect 248840 3544 248846 3556
rect 249886 3516 249892 3528
rect 248386 3488 249892 3516
rect 249886 3476 249892 3488
rect 249944 3476 249950 3528
rect 249978 3476 249984 3528
rect 250036 3516 250042 3528
rect 251082 3516 251088 3528
rect 250036 3488 251088 3516
rect 250036 3476 250042 3488
rect 251082 3476 251088 3488
rect 251140 3476 251146 3528
rect 251192 3516 251220 3556
rect 255866 3544 255872 3596
rect 255924 3584 255930 3596
rect 357434 3584 357440 3596
rect 255924 3556 357440 3584
rect 255924 3544 255930 3556
rect 357434 3544 357440 3556
rect 357492 3544 357498 3596
rect 362218 3584 362224 3596
rect 357544 3556 362224 3584
rect 353478 3516 353484 3528
rect 251192 3488 353484 3516
rect 353478 3476 353484 3488
rect 353536 3476 353542 3528
rect 354030 3476 354036 3528
rect 354088 3516 354094 3528
rect 354582 3516 354588 3528
rect 354088 3488 354588 3516
rect 354088 3476 354094 3488
rect 354582 3476 354588 3488
rect 354640 3476 354646 3528
rect 355137 3519 355195 3525
rect 355137 3485 355149 3519
rect 355183 3516 355195 3519
rect 357544 3516 357572 3556
rect 362218 3544 362224 3556
rect 362276 3544 362282 3596
rect 362310 3544 362316 3596
rect 362368 3584 362374 3596
rect 430574 3584 430580 3596
rect 362368 3556 430580 3584
rect 362368 3544 362374 3556
rect 430574 3544 430580 3556
rect 430632 3544 430638 3596
rect 430850 3544 430856 3596
rect 430908 3584 430914 3596
rect 432598 3584 432604 3596
rect 430908 3556 432604 3584
rect 430908 3544 430914 3556
rect 432598 3544 432604 3556
rect 432656 3544 432662 3596
rect 355183 3488 357572 3516
rect 355183 3485 355195 3488
rect 355137 3479 355195 3485
rect 361114 3476 361120 3528
rect 361172 3516 361178 3528
rect 363598 3516 363604 3528
rect 361172 3488 363604 3516
rect 361172 3476 361178 3488
rect 363598 3476 363604 3488
rect 363656 3476 363662 3528
rect 363693 3519 363751 3525
rect 363693 3485 363705 3519
rect 363739 3516 363751 3519
rect 422297 3519 422355 3525
rect 422297 3516 422309 3519
rect 363739 3488 422309 3516
rect 363739 3485 363751 3488
rect 363693 3479 363751 3485
rect 422297 3485 422309 3488
rect 422343 3485 422355 3519
rect 422297 3479 422355 3485
rect 422570 3476 422576 3528
rect 422628 3516 422634 3528
rect 423582 3516 423588 3528
rect 422628 3488 423588 3516
rect 422628 3476 422634 3488
rect 423582 3476 423588 3488
rect 423640 3476 423646 3528
rect 423766 3476 423772 3528
rect 423824 3516 423830 3528
rect 425698 3516 425704 3528
rect 423824 3488 425704 3516
rect 423824 3476 423830 3488
rect 425698 3476 425704 3488
rect 425756 3476 425762 3528
rect 427262 3476 427268 3528
rect 427320 3516 427326 3528
rect 428458 3516 428464 3528
rect 427320 3488 428464 3516
rect 427320 3476 427326 3488
rect 428458 3476 428464 3488
rect 428516 3476 428522 3528
rect 429654 3476 429660 3528
rect 429712 3516 429718 3528
rect 430482 3516 430488 3528
rect 429712 3488 430488 3516
rect 429712 3476 429718 3488
rect 430482 3476 430488 3488
rect 430540 3476 430546 3528
rect 432984 3516 433012 3624
rect 433076 3584 433104 3692
rect 436097 3689 436109 3723
rect 436143 3720 436155 3723
rect 440234 3720 440240 3732
rect 436143 3692 440240 3720
rect 436143 3689 436155 3692
rect 436097 3683 436155 3689
rect 440234 3680 440240 3692
rect 440292 3680 440298 3732
rect 433242 3612 433248 3664
rect 433300 3652 433306 3664
rect 433300 3624 439636 3652
rect 433300 3612 433306 3624
rect 436097 3587 436155 3593
rect 436097 3584 436109 3587
rect 433076 3556 436109 3584
rect 436097 3553 436109 3556
rect 436143 3553 436155 3587
rect 436097 3547 436155 3553
rect 437934 3544 437940 3596
rect 437992 3584 437998 3596
rect 439498 3584 439504 3596
rect 437992 3556 439504 3584
rect 437992 3544 437998 3556
rect 439498 3544 439504 3556
rect 439556 3544 439562 3596
rect 435358 3516 435364 3528
rect 432984 3488 435364 3516
rect 435358 3476 435364 3488
rect 435416 3476 435422 3528
rect 435542 3476 435548 3528
rect 435600 3516 435606 3528
rect 436002 3516 436008 3528
rect 435600 3488 436008 3516
rect 435600 3476 435606 3488
rect 436002 3476 436008 3488
rect 436060 3476 436066 3528
rect 436738 3476 436744 3528
rect 436796 3516 436802 3528
rect 438118 3516 438124 3528
rect 436796 3488 438124 3516
rect 436796 3476 436802 3488
rect 438118 3476 438124 3488
rect 438176 3476 438182 3528
rect 439608 3516 439636 3624
rect 440344 3584 440372 3760
rect 441522 3748 441528 3800
rect 441580 3788 441586 3800
rect 444929 3791 444987 3797
rect 444929 3788 444941 3791
rect 441580 3760 444941 3788
rect 441580 3748 441586 3760
rect 444929 3757 444941 3760
rect 444975 3757 444987 3791
rect 444929 3751 444987 3757
rect 445018 3748 445024 3800
rect 445076 3788 445082 3800
rect 447778 3788 447784 3800
rect 445076 3760 447784 3788
rect 445076 3748 445082 3760
rect 447778 3748 447784 3760
rect 447836 3748 447842 3800
rect 465718 3788 465724 3800
rect 451246 3760 465724 3788
rect 446214 3680 446220 3732
rect 446272 3720 446278 3732
rect 447042 3720 447048 3732
rect 446272 3692 447048 3720
rect 446272 3680 446278 3692
rect 447042 3680 447048 3692
rect 447100 3680 447106 3732
rect 447410 3680 447416 3732
rect 447468 3720 447474 3732
rect 451246 3720 451274 3760
rect 465718 3748 465724 3760
rect 465776 3748 465782 3800
rect 472250 3748 472256 3800
rect 472308 3788 472314 3800
rect 504358 3788 504364 3800
rect 472308 3760 504364 3788
rect 472308 3748 472314 3760
rect 504358 3748 504364 3760
rect 504416 3748 504422 3800
rect 509973 3791 510031 3797
rect 509973 3757 509985 3791
rect 510019 3788 510031 3791
rect 518158 3788 518164 3800
rect 510019 3760 518164 3788
rect 510019 3757 510031 3760
rect 509973 3751 510031 3757
rect 518158 3748 518164 3760
rect 518216 3748 518222 3800
rect 521838 3748 521844 3800
rect 521896 3788 521902 3800
rect 533338 3788 533344 3800
rect 521896 3760 533344 3788
rect 521896 3748 521902 3760
rect 533338 3748 533344 3760
rect 533396 3748 533402 3800
rect 447468 3692 451274 3720
rect 452013 3723 452071 3729
rect 447468 3680 447474 3692
rect 452013 3689 452025 3723
rect 452059 3720 452071 3723
rect 456058 3720 456064 3732
rect 452059 3692 456064 3720
rect 452059 3689 452071 3692
rect 452013 3683 452071 3689
rect 456058 3680 456064 3692
rect 456116 3680 456122 3732
rect 456886 3680 456892 3732
rect 456944 3720 456950 3732
rect 493318 3720 493324 3732
rect 456944 3692 493324 3720
rect 456944 3680 456950 3692
rect 493318 3680 493324 3692
rect 493376 3680 493382 3732
rect 499390 3680 499396 3732
rect 499448 3720 499454 3732
rect 502978 3720 502984 3732
rect 499448 3692 502984 3720
rect 499448 3680 499454 3692
rect 502978 3680 502984 3692
rect 503036 3680 503042 3732
rect 507670 3680 507676 3732
rect 507728 3720 507734 3732
rect 529290 3720 529296 3732
rect 507728 3692 529296 3720
rect 507728 3680 507734 3692
rect 529290 3680 529296 3692
rect 529348 3680 529354 3732
rect 536190 3720 536196 3732
rect 529952 3692 536196 3720
rect 440418 3612 440424 3664
rect 440476 3652 440482 3664
rect 479518 3652 479524 3664
rect 440476 3624 479524 3652
rect 440476 3612 440482 3624
rect 479518 3612 479524 3624
rect 479576 3612 479582 3664
rect 492306 3612 492312 3664
rect 492364 3652 492370 3664
rect 492364 3624 496860 3652
rect 492364 3612 492370 3624
rect 473998 3584 474004 3596
rect 440344 3556 474004 3584
rect 473998 3544 474004 3556
rect 474056 3544 474062 3596
rect 480441 3587 480499 3593
rect 480441 3553 480453 3587
rect 480487 3584 480499 3587
rect 487798 3584 487804 3596
rect 480487 3556 487804 3584
rect 480487 3553 480499 3556
rect 480441 3547 480499 3553
rect 487798 3544 487804 3556
rect 487856 3544 487862 3596
rect 488810 3544 488816 3596
rect 488868 3584 488874 3596
rect 489822 3584 489828 3596
rect 488868 3556 489828 3584
rect 488868 3544 488874 3556
rect 489822 3544 489828 3556
rect 489880 3544 489886 3596
rect 489914 3544 489920 3596
rect 489972 3584 489978 3596
rect 491202 3584 491208 3596
rect 489972 3556 491208 3584
rect 489972 3544 489978 3556
rect 491202 3544 491208 3556
rect 491260 3544 491266 3596
rect 493502 3544 493508 3596
rect 493560 3584 493566 3596
rect 493962 3584 493968 3596
rect 493560 3556 493968 3584
rect 493560 3544 493566 3556
rect 493962 3544 493968 3556
rect 494020 3544 494026 3596
rect 495894 3544 495900 3596
rect 495952 3584 495958 3596
rect 496722 3584 496728 3596
rect 495952 3556 496728 3584
rect 495952 3544 495958 3556
rect 496722 3544 496728 3556
rect 496780 3544 496786 3596
rect 496832 3584 496860 3624
rect 498194 3612 498200 3664
rect 498252 3652 498258 3664
rect 522390 3652 522396 3664
rect 498252 3624 522396 3652
rect 498252 3612 498258 3624
rect 522390 3612 522396 3624
rect 522448 3612 522454 3664
rect 529952 3652 529980 3692
rect 536190 3680 536196 3692
rect 536248 3680 536254 3732
rect 546678 3680 546684 3732
rect 546736 3720 546742 3732
rect 548518 3720 548524 3732
rect 546736 3692 548524 3720
rect 546736 3680 546742 3692
rect 548518 3680 548524 3692
rect 548576 3680 548582 3732
rect 528526 3624 529980 3652
rect 509973 3587 510031 3593
rect 509973 3584 509985 3587
rect 496832 3556 509985 3584
rect 509973 3553 509985 3556
rect 510019 3553 510031 3587
rect 509973 3547 510031 3553
rect 510062 3544 510068 3596
rect 510120 3584 510126 3596
rect 525058 3584 525064 3596
rect 510120 3556 525064 3584
rect 510120 3544 510126 3556
rect 525058 3544 525064 3556
rect 525116 3544 525122 3596
rect 525426 3544 525432 3596
rect 525484 3584 525490 3596
rect 528526 3584 528554 3624
rect 543182 3612 543188 3664
rect 543240 3652 543246 3664
rect 544378 3652 544384 3664
rect 543240 3624 544384 3652
rect 543240 3612 543246 3624
rect 544378 3612 544384 3624
rect 544436 3612 544442 3664
rect 536098 3584 536104 3596
rect 525484 3556 528554 3584
rect 530136 3556 536104 3584
rect 525484 3544 525490 3556
rect 470965 3519 471023 3525
rect 470965 3516 470977 3519
rect 439608 3488 470977 3516
rect 470965 3485 470977 3488
rect 471011 3485 471023 3519
rect 470965 3479 471023 3485
rect 471054 3476 471060 3528
rect 471112 3516 471118 3528
rect 478046 3516 478052 3528
rect 471112 3488 478052 3516
rect 471112 3476 471118 3488
rect 478046 3476 478052 3488
rect 478104 3476 478110 3528
rect 479334 3476 479340 3528
rect 479392 3516 479398 3528
rect 480162 3516 480168 3528
rect 479392 3488 480168 3516
rect 479392 3476 479398 3488
rect 480162 3476 480168 3488
rect 480220 3476 480226 3528
rect 482830 3476 482836 3528
rect 482888 3516 482894 3528
rect 482888 3488 483060 3516
rect 482888 3476 482894 3488
rect 186406 3448 186412 3460
rect 10008 3352 14596 3380
rect 14660 3420 186412 3448
rect 10008 3340 10014 3352
rect 14660 3312 14688 3420
rect 186406 3408 186412 3420
rect 186464 3408 186470 3460
rect 189718 3408 189724 3460
rect 189776 3448 189782 3460
rect 190362 3448 190368 3460
rect 189776 3420 190368 3448
rect 189776 3408 189782 3420
rect 190362 3408 190368 3420
rect 190420 3408 190426 3460
rect 199102 3408 199108 3460
rect 199160 3448 199166 3460
rect 200022 3448 200028 3460
rect 199160 3420 200028 3448
rect 199160 3408 199166 3420
rect 200022 3408 200028 3420
rect 200080 3408 200086 3460
rect 200298 3408 200304 3460
rect 200356 3448 200362 3460
rect 230937 3451 230995 3457
rect 230937 3448 230949 3451
rect 200356 3420 230949 3448
rect 200356 3408 200362 3420
rect 230937 3417 230949 3420
rect 230983 3417 230995 3451
rect 230937 3411 230995 3417
rect 231026 3408 231032 3460
rect 231084 3448 231090 3460
rect 231762 3448 231768 3460
rect 231084 3420 231768 3448
rect 231084 3408 231090 3420
rect 231762 3408 231768 3420
rect 231820 3408 231826 3460
rect 232222 3408 232228 3460
rect 232280 3448 232286 3460
rect 241609 3451 241667 3457
rect 241609 3448 241621 3451
rect 232280 3420 241621 3448
rect 232280 3408 232286 3420
rect 241609 3417 241621 3420
rect 241655 3417 241667 3451
rect 241609 3411 241667 3417
rect 241698 3408 241704 3460
rect 241756 3448 241762 3460
rect 340049 3451 340107 3457
rect 340049 3448 340061 3451
rect 241756 3420 340061 3448
rect 241756 3408 241762 3420
rect 340049 3417 340061 3420
rect 340095 3417 340107 3451
rect 340049 3411 340107 3417
rect 344554 3408 344560 3460
rect 344612 3448 344618 3460
rect 345658 3448 345664 3460
rect 344612 3420 345664 3448
rect 344612 3408 344618 3420
rect 345658 3408 345664 3420
rect 345716 3408 345722 3460
rect 348050 3408 348056 3460
rect 348108 3448 348114 3460
rect 413005 3451 413063 3457
rect 413005 3448 413017 3451
rect 348108 3420 413017 3448
rect 348108 3408 348114 3420
rect 413005 3417 413017 3420
rect 413051 3417 413063 3451
rect 413005 3411 413063 3417
rect 413094 3408 413100 3460
rect 413152 3448 413158 3460
rect 414658 3448 414664 3460
rect 413152 3420 414664 3448
rect 413152 3408 413158 3420
rect 414658 3408 414664 3420
rect 414716 3408 414722 3460
rect 415486 3408 415492 3460
rect 415544 3448 415550 3460
rect 416682 3448 416688 3460
rect 415544 3420 416688 3448
rect 415544 3408 415550 3420
rect 416682 3408 416688 3420
rect 416740 3408 416746 3460
rect 421374 3408 421380 3460
rect 421432 3448 421438 3460
rect 424318 3448 424324 3460
rect 421432 3420 424324 3448
rect 421432 3408 421438 3420
rect 424318 3408 424324 3420
rect 424376 3408 424382 3460
rect 426158 3408 426164 3460
rect 426216 3448 426222 3460
rect 474734 3448 474740 3460
rect 426216 3420 474740 3448
rect 426216 3408 426222 3420
rect 474734 3408 474740 3420
rect 474792 3408 474798 3460
rect 478230 3448 478236 3460
rect 474844 3420 478236 3448
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 17218 3380 17224 3392
rect 15988 3352 17224 3380
rect 15988 3340 15994 3352
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 32398 3340 32404 3392
rect 32456 3380 32462 3392
rect 33778 3380 33784 3392
rect 32456 3352 33784 3380
rect 32456 3340 32462 3352
rect 33778 3340 33784 3352
rect 33836 3340 33842 3392
rect 39574 3340 39580 3392
rect 39632 3380 39638 3392
rect 43438 3380 43444 3392
rect 39632 3352 43444 3380
rect 39632 3340 39638 3352
rect 43438 3340 43444 3352
rect 43496 3340 43502 3392
rect 45462 3340 45468 3392
rect 45520 3380 45526 3392
rect 54478 3380 54484 3392
rect 45520 3352 54484 3380
rect 45520 3340 45526 3352
rect 54478 3340 54484 3352
rect 54536 3340 54542 3392
rect 74994 3340 75000 3392
rect 75052 3380 75058 3392
rect 214558 3380 214564 3392
rect 75052 3352 214564 3380
rect 75052 3340 75058 3352
rect 214558 3340 214564 3352
rect 214616 3340 214622 3392
rect 222746 3340 222752 3392
rect 222804 3380 222810 3392
rect 223482 3380 223488 3392
rect 222804 3352 223488 3380
rect 222804 3340 222810 3352
rect 223482 3340 223488 3352
rect 223540 3340 223546 3392
rect 238110 3340 238116 3392
rect 238168 3380 238174 3392
rect 249058 3380 249064 3392
rect 238168 3352 249064 3380
rect 238168 3340 238174 3352
rect 249058 3340 249064 3352
rect 249116 3340 249122 3392
rect 252370 3340 252376 3392
rect 252428 3380 252434 3392
rect 278038 3380 278044 3392
rect 252428 3352 278044 3380
rect 252428 3340 252434 3352
rect 278038 3340 278044 3352
rect 278096 3340 278102 3392
rect 278314 3340 278320 3392
rect 278372 3380 278378 3392
rect 280798 3380 280804 3392
rect 278372 3352 280804 3380
rect 278372 3340 278378 3352
rect 280798 3340 280804 3352
rect 280856 3340 280862 3392
rect 283098 3340 283104 3392
rect 283156 3380 283162 3392
rect 286318 3380 286324 3392
rect 283156 3352 286324 3380
rect 283156 3340 283162 3352
rect 286318 3340 286324 3352
rect 286376 3340 286382 3392
rect 286594 3340 286600 3392
rect 286652 3380 286658 3392
rect 320818 3380 320824 3392
rect 286652 3352 320824 3380
rect 286652 3340 286658 3352
rect 320818 3340 320824 3352
rect 320876 3340 320882 3392
rect 322106 3340 322112 3392
rect 322164 3380 322170 3392
rect 323578 3380 323584 3392
rect 322164 3352 323584 3380
rect 322164 3340 322170 3352
rect 323578 3340 323584 3352
rect 323636 3340 323642 3392
rect 330386 3340 330392 3392
rect 330444 3380 330450 3392
rect 331858 3380 331864 3392
rect 330444 3352 331864 3380
rect 330444 3340 330450 3352
rect 331858 3340 331864 3352
rect 331916 3340 331922 3392
rect 331968 3352 404676 3380
rect 9876 3284 14688 3312
rect 41874 3272 41880 3324
rect 41932 3312 41938 3324
rect 50065 3315 50123 3321
rect 50065 3312 50077 3315
rect 41932 3284 50077 3312
rect 41932 3272 41938 3284
rect 50065 3281 50077 3284
rect 50111 3281 50123 3315
rect 50065 3275 50123 3281
rect 50154 3272 50160 3324
rect 50212 3312 50218 3324
rect 79318 3312 79324 3324
rect 50212 3284 79324 3312
rect 50212 3272 50218 3284
rect 79318 3272 79324 3284
rect 79376 3272 79382 3324
rect 80882 3272 80888 3324
rect 80940 3312 80946 3324
rect 81342 3312 81348 3324
rect 80940 3284 81348 3312
rect 80940 3272 80946 3284
rect 81342 3272 81348 3284
rect 81400 3272 81406 3324
rect 84470 3272 84476 3324
rect 84528 3312 84534 3324
rect 86218 3312 86224 3324
rect 84528 3284 86224 3312
rect 84528 3272 84534 3284
rect 86218 3272 86224 3284
rect 86276 3272 86282 3324
rect 87966 3272 87972 3324
rect 88024 3312 88030 3324
rect 88978 3312 88984 3324
rect 88024 3284 88984 3312
rect 88024 3272 88030 3284
rect 88978 3272 88984 3284
rect 89036 3272 89042 3324
rect 89162 3272 89168 3324
rect 89220 3312 89226 3324
rect 90358 3312 90364 3324
rect 89220 3284 90364 3312
rect 89220 3272 89226 3284
rect 90358 3272 90364 3284
rect 90416 3272 90422 3324
rect 91554 3272 91560 3324
rect 91612 3312 91618 3324
rect 93118 3312 93124 3324
rect 91612 3284 93124 3312
rect 91612 3272 91618 3284
rect 93118 3272 93124 3284
rect 93176 3272 93182 3324
rect 93213 3315 93271 3321
rect 93213 3281 93225 3315
rect 93259 3312 93271 3315
rect 217318 3312 217324 3324
rect 93259 3284 217324 3312
rect 93259 3281 93271 3284
rect 93213 3275 93271 3281
rect 217318 3272 217324 3284
rect 217376 3272 217382 3324
rect 228726 3272 228732 3324
rect 228784 3312 228790 3324
rect 238018 3312 238024 3324
rect 228784 3284 238024 3312
rect 228784 3272 228790 3284
rect 238018 3272 238024 3284
rect 238076 3272 238082 3324
rect 242158 3312 242164 3324
rect 238726 3284 242164 3312
rect 18230 3204 18236 3256
rect 18288 3244 18294 3256
rect 22738 3244 22744 3256
rect 18288 3216 22744 3244
rect 18288 3204 18294 3216
rect 22738 3204 22744 3216
rect 22796 3204 22802 3256
rect 23014 3204 23020 3256
rect 23072 3244 23078 3256
rect 25498 3244 25504 3256
rect 23072 3216 25504 3244
rect 23072 3204 23078 3216
rect 25498 3204 25504 3216
rect 25556 3204 25562 3256
rect 57238 3204 57244 3256
rect 57296 3244 57302 3256
rect 83458 3244 83464 3256
rect 57296 3216 83464 3244
rect 57296 3204 57302 3216
rect 83458 3204 83464 3216
rect 83516 3204 83522 3256
rect 85666 3204 85672 3256
rect 85724 3244 85730 3256
rect 220078 3244 220084 3256
rect 85724 3216 220084 3244
rect 85724 3204 85730 3216
rect 220078 3204 220084 3216
rect 220136 3204 220142 3256
rect 235810 3204 235816 3256
rect 235868 3244 235874 3256
rect 238726 3244 238754 3284
rect 242158 3272 242164 3284
rect 242216 3272 242222 3324
rect 246390 3272 246396 3324
rect 246448 3312 246454 3324
rect 269850 3312 269856 3324
rect 246448 3284 269856 3312
rect 246448 3272 246454 3284
rect 269850 3272 269856 3284
rect 269908 3272 269914 3324
rect 274818 3272 274824 3324
rect 274876 3312 274882 3324
rect 276750 3312 276756 3324
rect 274876 3284 276756 3312
rect 274876 3272 274882 3284
rect 276750 3272 276756 3284
rect 276808 3272 276814 3324
rect 279421 3315 279479 3321
rect 279421 3281 279433 3315
rect 279467 3312 279479 3315
rect 287698 3312 287704 3324
rect 279467 3284 287704 3312
rect 279467 3281 279479 3284
rect 279421 3275 279479 3281
rect 287698 3272 287704 3284
rect 287756 3272 287762 3324
rect 290182 3272 290188 3324
rect 290240 3312 290246 3324
rect 309778 3312 309784 3324
rect 290240 3284 309784 3312
rect 290240 3272 290246 3284
rect 309778 3272 309784 3284
rect 309836 3272 309842 3324
rect 311434 3272 311440 3324
rect 311492 3312 311498 3324
rect 312630 3312 312636 3324
rect 311492 3284 312636 3312
rect 311492 3272 311498 3284
rect 312630 3272 312636 3284
rect 312688 3272 312694 3324
rect 312722 3272 312728 3324
rect 312780 3312 312786 3324
rect 325697 3315 325755 3321
rect 325697 3312 325709 3315
rect 312780 3284 325709 3312
rect 312780 3272 312786 3284
rect 325697 3281 325709 3284
rect 325743 3281 325755 3315
rect 325697 3275 325755 3281
rect 326798 3272 326804 3324
rect 326856 3312 326862 3324
rect 331968 3312 331996 3352
rect 388073 3315 388131 3321
rect 388073 3312 388085 3315
rect 326856 3284 331996 3312
rect 335326 3284 388085 3312
rect 326856 3272 326862 3284
rect 240962 3244 240968 3256
rect 235868 3216 238754 3244
rect 239232 3216 240968 3244
rect 235868 3204 235874 3216
rect 64322 3136 64328 3188
rect 64380 3176 64386 3188
rect 87598 3176 87604 3188
rect 64380 3148 87604 3176
rect 64380 3136 64386 3148
rect 87598 3136 87604 3148
rect 87656 3136 87662 3188
rect 92750 3136 92756 3188
rect 92808 3176 92814 3188
rect 221458 3176 221464 3188
rect 92808 3148 221464 3176
rect 92808 3136 92814 3148
rect 221458 3136 221464 3148
rect 221516 3136 221522 3188
rect 230937 3179 230995 3185
rect 230937 3145 230949 3179
rect 230983 3176 230995 3179
rect 239232 3176 239260 3216
rect 240962 3204 240968 3216
rect 241020 3204 241026 3256
rect 242894 3204 242900 3256
rect 242952 3244 242958 3256
rect 260098 3244 260104 3256
rect 242952 3216 260104 3244
rect 242952 3204 242958 3216
rect 260098 3204 260104 3216
rect 260156 3204 260162 3256
rect 260650 3204 260656 3256
rect 260708 3244 260714 3256
rect 268470 3244 268476 3256
rect 260708 3216 268476 3244
rect 260708 3204 260714 3216
rect 268470 3204 268476 3216
rect 268528 3204 268534 3256
rect 273622 3204 273628 3256
rect 273680 3244 273686 3256
rect 282178 3244 282184 3256
rect 273680 3216 282184 3244
rect 273680 3204 273686 3216
rect 282178 3204 282184 3216
rect 282236 3204 282242 3256
rect 291378 3204 291384 3256
rect 291436 3244 291442 3256
rect 297177 3247 297235 3253
rect 297177 3244 297189 3247
rect 291436 3216 297189 3244
rect 291436 3204 291442 3216
rect 297177 3213 297189 3216
rect 297223 3213 297235 3247
rect 297177 3207 297235 3213
rect 297266 3204 297272 3256
rect 297324 3244 297330 3256
rect 304258 3244 304264 3256
rect 297324 3216 304264 3244
rect 297324 3204 297330 3216
rect 304258 3204 304264 3216
rect 304316 3204 304322 3256
rect 304350 3204 304356 3256
rect 304408 3244 304414 3256
rect 305730 3244 305736 3256
rect 304408 3216 305736 3244
rect 304408 3204 304414 3216
rect 305730 3204 305736 3216
rect 305788 3204 305794 3256
rect 316129 3247 316187 3253
rect 316129 3244 316141 3247
rect 305932 3216 316141 3244
rect 230983 3148 239260 3176
rect 230983 3145 230995 3148
rect 230937 3139 230995 3145
rect 239306 3136 239312 3188
rect 239364 3176 239370 3188
rect 244918 3176 244924 3188
rect 239364 3148 244924 3176
rect 239364 3136 239370 3148
rect 244918 3136 244924 3148
rect 244976 3136 244982 3188
rect 245194 3136 245200 3188
rect 245252 3176 245258 3188
rect 255958 3176 255964 3188
rect 245252 3148 255964 3176
rect 245252 3136 245258 3148
rect 255958 3136 255964 3148
rect 256016 3136 256022 3188
rect 258077 3179 258135 3185
rect 258077 3145 258089 3179
rect 258123 3176 258135 3179
rect 266998 3176 267004 3188
rect 258123 3148 267004 3176
rect 258123 3145 258135 3148
rect 258077 3139 258135 3145
rect 266998 3136 267004 3148
rect 267056 3136 267062 3188
rect 294874 3136 294880 3188
rect 294932 3176 294938 3188
rect 294932 3148 301544 3176
rect 294932 3136 294938 3148
rect 71498 3068 71504 3120
rect 71556 3108 71562 3120
rect 98546 3108 98552 3120
rect 71556 3080 98552 3108
rect 71556 3068 71562 3080
rect 98546 3068 98552 3080
rect 98604 3068 98610 3120
rect 98638 3068 98644 3120
rect 98696 3108 98702 3120
rect 99282 3108 99288 3120
rect 98696 3080 99288 3108
rect 98696 3068 98702 3080
rect 99282 3068 99288 3080
rect 99340 3068 99346 3120
rect 102226 3068 102232 3120
rect 102284 3108 102290 3120
rect 104158 3108 104164 3120
rect 102284 3080 104164 3108
rect 102284 3068 102290 3080
rect 104158 3068 104164 3080
rect 104216 3068 104222 3120
rect 106918 3068 106924 3120
rect 106976 3108 106982 3120
rect 107562 3108 107568 3120
rect 106976 3080 107568 3108
rect 106976 3068 106982 3080
rect 107562 3068 107568 3080
rect 107620 3068 107626 3120
rect 109310 3068 109316 3120
rect 109368 3108 109374 3120
rect 111058 3108 111064 3120
rect 109368 3080 111064 3108
rect 109368 3068 109374 3080
rect 111058 3068 111064 3080
rect 111116 3068 111122 3120
rect 224218 3108 224224 3120
rect 111168 3080 224224 3108
rect 46658 3000 46664 3052
rect 46716 3040 46722 3052
rect 50338 3040 50344 3052
rect 46716 3012 50344 3040
rect 46716 3000 46722 3012
rect 50338 3000 50344 3012
rect 50396 3000 50402 3052
rect 78582 3000 78588 3052
rect 78640 3040 78646 3052
rect 78640 3012 93854 3040
rect 78640 3000 78646 3012
rect 82078 2932 82084 2984
rect 82136 2972 82142 2984
rect 93213 2975 93271 2981
rect 93213 2972 93225 2975
rect 82136 2944 93225 2972
rect 82136 2932 82142 2944
rect 93213 2941 93225 2944
rect 93259 2941 93271 2975
rect 93213 2935 93271 2941
rect 93826 2904 93854 3012
rect 99834 3000 99840 3052
rect 99892 3040 99898 3052
rect 111168 3040 111196 3080
rect 224218 3068 224224 3080
rect 224276 3068 224282 3120
rect 268838 3068 268844 3120
rect 268896 3108 268902 3120
rect 276658 3108 276664 3120
rect 268896 3080 276664 3108
rect 268896 3068 268902 3080
rect 276658 3068 276664 3080
rect 276716 3068 276722 3120
rect 280706 3068 280712 3120
rect 280764 3108 280770 3120
rect 284938 3108 284944 3120
rect 280764 3080 284944 3108
rect 280764 3068 280770 3080
rect 284938 3068 284944 3080
rect 284996 3068 285002 3120
rect 287790 3068 287796 3120
rect 287848 3108 287854 3120
rect 295978 3108 295984 3120
rect 287848 3080 295984 3108
rect 287848 3068 287854 3080
rect 295978 3068 295984 3080
rect 296036 3068 296042 3120
rect 226978 3040 226984 3052
rect 99892 3012 111196 3040
rect 113146 3012 226984 3040
rect 99892 3000 99898 3012
rect 96246 2932 96252 2984
rect 96304 2972 96310 2984
rect 101398 2972 101404 2984
rect 96304 2944 101404 2972
rect 96304 2932 96310 2944
rect 101398 2932 101404 2944
rect 101456 2932 101462 2984
rect 105722 2932 105728 2984
rect 105780 2972 105786 2984
rect 108298 2972 108304 2984
rect 105780 2944 108304 2972
rect 105780 2932 105786 2944
rect 108298 2932 108304 2944
rect 108356 2932 108362 2984
rect 110506 2932 110512 2984
rect 110564 2972 110570 2984
rect 113146 2972 113174 3012
rect 226978 3000 226984 3012
rect 227036 3000 227042 3052
rect 296070 3000 296076 3052
rect 296128 3040 296134 3052
rect 296622 3040 296628 3052
rect 296128 3012 296628 3040
rect 296128 3000 296134 3012
rect 296622 3000 296628 3012
rect 296680 3000 296686 3052
rect 301516 3040 301544 3148
rect 301958 3068 301964 3120
rect 302016 3108 302022 3120
rect 305932 3108 305960 3216
rect 316129 3213 316141 3216
rect 316175 3213 316187 3247
rect 316129 3207 316187 3213
rect 316218 3204 316224 3256
rect 316276 3244 316282 3256
rect 322198 3244 322204 3256
rect 316276 3216 322204 3244
rect 316276 3204 316282 3216
rect 322198 3204 322204 3216
rect 322256 3204 322262 3256
rect 323302 3204 323308 3256
rect 323360 3244 323366 3256
rect 327718 3244 327724 3256
rect 323360 3216 327724 3244
rect 323360 3204 323366 3216
rect 327718 3204 327724 3216
rect 327776 3204 327782 3256
rect 332045 3247 332103 3253
rect 332045 3213 332057 3247
rect 332091 3244 332103 3247
rect 335326 3244 335354 3284
rect 388073 3281 388085 3284
rect 388119 3281 388131 3315
rect 388073 3275 388131 3281
rect 391842 3272 391848 3324
rect 391900 3312 391906 3324
rect 392670 3312 392676 3324
rect 391900 3284 392676 3312
rect 391900 3272 391906 3284
rect 392670 3272 392676 3284
rect 392728 3272 392734 3324
rect 395338 3272 395344 3324
rect 395396 3312 395402 3324
rect 395982 3312 395988 3324
rect 395396 3284 395988 3312
rect 395396 3272 395402 3284
rect 395982 3272 395988 3284
rect 396040 3272 396046 3324
rect 398926 3272 398932 3324
rect 398984 3312 398990 3324
rect 400858 3312 400864 3324
rect 398984 3284 400864 3312
rect 398984 3272 398990 3284
rect 400858 3272 400864 3284
rect 400916 3272 400922 3324
rect 401318 3272 401324 3324
rect 401376 3312 401382 3324
rect 402238 3312 402244 3324
rect 401376 3284 402244 3312
rect 401376 3272 401382 3284
rect 402238 3272 402244 3284
rect 402296 3272 402302 3324
rect 402333 3315 402391 3321
rect 402333 3281 402345 3315
rect 402379 3312 402391 3315
rect 404081 3315 404139 3321
rect 404081 3312 404093 3315
rect 402379 3284 404093 3312
rect 402379 3281 402391 3284
rect 402333 3275 402391 3281
rect 404081 3281 404093 3284
rect 404127 3281 404139 3315
rect 404081 3275 404139 3281
rect 332091 3216 335354 3244
rect 339865 3247 339923 3253
rect 332091 3213 332103 3216
rect 332045 3207 332103 3213
rect 339865 3213 339877 3247
rect 339911 3244 339923 3247
rect 404541 3247 404599 3253
rect 404541 3244 404553 3247
rect 339911 3216 404553 3244
rect 339911 3213 339923 3216
rect 339865 3207 339923 3213
rect 404541 3213 404553 3216
rect 404587 3213 404599 3247
rect 404648 3244 404676 3352
rect 406010 3340 406016 3392
rect 406068 3380 406074 3392
rect 407022 3380 407028 3392
rect 406068 3352 407028 3380
rect 406068 3340 406074 3352
rect 407022 3340 407028 3352
rect 407080 3340 407086 3392
rect 407206 3340 407212 3392
rect 407264 3380 407270 3392
rect 411898 3380 411904 3392
rect 407264 3352 411904 3380
rect 407264 3340 407270 3352
rect 411898 3340 411904 3352
rect 411956 3340 411962 3392
rect 414290 3340 414296 3392
rect 414348 3380 414354 3392
rect 416038 3380 416044 3392
rect 414348 3352 416044 3380
rect 414348 3340 414354 3352
rect 416038 3340 416044 3352
rect 416096 3340 416102 3392
rect 422941 3383 422999 3389
rect 422941 3349 422953 3383
rect 422987 3380 422999 3383
rect 422987 3352 462728 3380
rect 422987 3349 422999 3352
rect 422941 3343 422999 3349
rect 404814 3272 404820 3324
rect 404872 3312 404878 3324
rect 452013 3315 452071 3321
rect 452013 3312 452025 3315
rect 404872 3284 452025 3312
rect 404872 3272 404878 3284
rect 452013 3281 452025 3284
rect 452059 3281 452071 3315
rect 452013 3275 452071 3281
rect 452102 3272 452108 3324
rect 452160 3312 452166 3324
rect 453298 3312 453304 3324
rect 452160 3284 453304 3312
rect 452160 3272 452166 3284
rect 453298 3272 453304 3284
rect 453356 3272 453362 3324
rect 455690 3272 455696 3324
rect 455748 3312 455754 3324
rect 457438 3312 457444 3324
rect 455748 3284 457444 3312
rect 455748 3272 455754 3284
rect 457438 3272 457444 3284
rect 457496 3272 457502 3324
rect 406378 3244 406384 3256
rect 404648 3216 406384 3244
rect 404541 3207 404599 3213
rect 406378 3204 406384 3216
rect 406436 3204 406442 3256
rect 410794 3204 410800 3256
rect 410852 3244 410858 3256
rect 416593 3247 416651 3253
rect 416593 3244 416605 3247
rect 410852 3216 416605 3244
rect 410852 3204 410858 3216
rect 416593 3213 416605 3216
rect 416639 3213 416651 3247
rect 416593 3207 416651 3213
rect 416682 3204 416688 3256
rect 416740 3244 416746 3256
rect 418798 3244 418804 3256
rect 416740 3216 418804 3244
rect 416740 3204 416746 3216
rect 418798 3204 418804 3216
rect 418856 3204 418862 3256
rect 418982 3204 418988 3256
rect 419040 3244 419046 3256
rect 462593 3247 462651 3253
rect 462593 3244 462605 3247
rect 419040 3216 462605 3244
rect 419040 3204 419046 3216
rect 462593 3213 462605 3216
rect 462639 3213 462651 3247
rect 462700 3244 462728 3352
rect 462774 3340 462780 3392
rect 462832 3380 462838 3392
rect 464338 3380 464344 3392
rect 462832 3352 464344 3380
rect 462832 3340 462838 3352
rect 464338 3340 464344 3352
rect 464396 3340 464402 3392
rect 465166 3340 465172 3392
rect 465224 3380 465230 3392
rect 466362 3380 466368 3392
rect 465224 3352 466368 3380
rect 465224 3340 465230 3352
rect 466362 3340 466368 3352
rect 466420 3340 466426 3392
rect 470965 3383 471023 3389
rect 470965 3349 470977 3383
rect 471011 3380 471023 3383
rect 474844 3380 474872 3420
rect 478230 3408 478236 3420
rect 478288 3408 478294 3460
rect 481726 3408 481732 3460
rect 481784 3448 481790 3460
rect 482922 3448 482928 3460
rect 481784 3420 482928 3448
rect 481784 3408 481790 3420
rect 482922 3408 482928 3420
rect 482980 3408 482986 3460
rect 483032 3448 483060 3488
rect 485222 3476 485228 3528
rect 485280 3516 485286 3528
rect 485682 3516 485688 3528
rect 485280 3488 485688 3516
rect 485280 3476 485286 3488
rect 485682 3476 485688 3488
rect 485740 3476 485746 3528
rect 487614 3476 487620 3528
rect 487672 3516 487678 3528
rect 489178 3516 489184 3528
rect 487672 3488 489184 3516
rect 487672 3476 487678 3488
rect 489178 3476 489184 3488
rect 489236 3476 489242 3528
rect 502889 3519 502947 3525
rect 502889 3516 502901 3519
rect 489288 3488 502901 3516
rect 489288 3448 489316 3488
rect 502889 3485 502901 3488
rect 502935 3485 502947 3519
rect 502889 3479 502947 3485
rect 502978 3476 502984 3528
rect 503036 3516 503042 3528
rect 503622 3516 503628 3528
rect 503036 3488 503628 3516
rect 503036 3476 503042 3488
rect 503622 3476 503628 3488
rect 503680 3476 503686 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507762 3516 507768 3528
rect 506532 3488 507768 3516
rect 506532 3476 506538 3488
rect 507762 3476 507768 3488
rect 507820 3476 507826 3528
rect 511258 3476 511264 3528
rect 511316 3516 511322 3528
rect 511902 3516 511908 3528
rect 511316 3488 511908 3516
rect 511316 3476 511322 3488
rect 511902 3476 511908 3488
rect 511960 3476 511966 3528
rect 512454 3476 512460 3528
rect 512512 3516 512518 3528
rect 513282 3516 513288 3528
rect 512512 3488 513288 3516
rect 512512 3476 512518 3488
rect 513282 3476 513288 3488
rect 513340 3476 513346 3528
rect 513558 3476 513564 3528
rect 513616 3516 513622 3528
rect 515398 3516 515404 3528
rect 513616 3488 515404 3516
rect 513616 3476 513622 3488
rect 515398 3476 515404 3488
rect 515456 3476 515462 3528
rect 518342 3476 518348 3528
rect 518400 3516 518406 3528
rect 518802 3516 518808 3528
rect 518400 3488 518808 3516
rect 518400 3476 518406 3488
rect 518802 3476 518808 3488
rect 518860 3476 518866 3528
rect 519538 3476 519544 3528
rect 519596 3516 519602 3528
rect 520182 3516 520188 3528
rect 519596 3488 520188 3516
rect 519596 3476 519602 3488
rect 520182 3476 520188 3488
rect 520240 3476 520246 3528
rect 520734 3476 520740 3528
rect 520792 3516 520798 3528
rect 521562 3516 521568 3528
rect 520792 3488 521568 3516
rect 520792 3476 520798 3488
rect 521562 3476 521568 3488
rect 521620 3476 521626 3528
rect 523034 3476 523040 3528
rect 523092 3516 523098 3528
rect 526438 3516 526444 3528
rect 523092 3488 526444 3516
rect 523092 3476 523098 3488
rect 526438 3476 526444 3488
rect 526496 3476 526502 3528
rect 526622 3476 526628 3528
rect 526680 3516 526686 3528
rect 527082 3516 527088 3528
rect 526680 3488 527088 3516
rect 526680 3476 526686 3488
rect 527082 3476 527088 3488
rect 527140 3476 527146 3528
rect 527818 3476 527824 3528
rect 527876 3516 527882 3528
rect 530136 3516 530164 3556
rect 536098 3544 536104 3556
rect 536156 3544 536162 3596
rect 549070 3544 549076 3596
rect 549128 3584 549134 3596
rect 554038 3584 554044 3596
rect 549128 3556 554044 3584
rect 549128 3544 549134 3556
rect 554038 3544 554044 3556
rect 554096 3544 554102 3596
rect 565630 3544 565636 3596
rect 565688 3584 565694 3596
rect 569310 3584 569316 3596
rect 565688 3556 569316 3584
rect 565688 3544 565694 3556
rect 569310 3544 569316 3556
rect 569368 3544 569374 3596
rect 527876 3488 530164 3516
rect 527876 3476 527882 3488
rect 534902 3476 534908 3528
rect 534960 3516 534966 3528
rect 535362 3516 535368 3528
rect 534960 3488 535368 3516
rect 534960 3476 534966 3488
rect 535362 3476 535368 3488
rect 535420 3476 535426 3528
rect 537202 3476 537208 3528
rect 537260 3516 537266 3528
rect 538122 3516 538128 3528
rect 537260 3488 538128 3516
rect 537260 3476 537266 3488
rect 538122 3476 538128 3488
rect 538180 3476 538186 3528
rect 538398 3476 538404 3528
rect 538456 3516 538462 3528
rect 539502 3516 539508 3528
rect 538456 3488 539508 3516
rect 538456 3476 538462 3488
rect 539502 3476 539508 3488
rect 539560 3476 539566 3528
rect 541986 3476 541992 3528
rect 542044 3516 542050 3528
rect 542998 3516 543004 3528
rect 542044 3488 543004 3516
rect 542044 3476 542050 3488
rect 542998 3476 543004 3488
rect 543056 3476 543062 3528
rect 544378 3476 544384 3528
rect 544436 3516 544442 3528
rect 545022 3516 545028 3528
rect 544436 3488 545028 3516
rect 544436 3476 544442 3488
rect 545022 3476 545028 3488
rect 545080 3476 545086 3528
rect 545482 3476 545488 3528
rect 545540 3516 545546 3528
rect 547138 3516 547144 3528
rect 545540 3488 547144 3516
rect 545540 3476 545546 3488
rect 547138 3476 547144 3488
rect 547196 3476 547202 3528
rect 547874 3476 547880 3528
rect 547932 3516 547938 3528
rect 549162 3516 549168 3528
rect 547932 3488 549168 3516
rect 547932 3476 547938 3488
rect 549162 3476 549168 3488
rect 549220 3476 549226 3528
rect 550266 3476 550272 3528
rect 550324 3516 550330 3528
rect 551278 3516 551284 3528
rect 550324 3488 551284 3516
rect 550324 3476 550330 3488
rect 551278 3476 551284 3488
rect 551336 3476 551342 3528
rect 551462 3476 551468 3528
rect 551520 3516 551526 3528
rect 551922 3516 551928 3528
rect 551520 3488 551928 3516
rect 551520 3476 551526 3488
rect 551922 3476 551928 3488
rect 551980 3476 551986 3528
rect 556154 3476 556160 3528
rect 556212 3516 556218 3528
rect 557442 3516 557448 3528
rect 556212 3488 557448 3516
rect 556212 3476 556218 3488
rect 557442 3476 557448 3488
rect 557500 3476 557506 3528
rect 560846 3476 560852 3528
rect 560904 3516 560910 3528
rect 561582 3516 561588 3528
rect 560904 3488 561588 3516
rect 560904 3476 560910 3488
rect 561582 3476 561588 3488
rect 561640 3476 561646 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565722 3516 565728 3528
rect 564492 3488 565728 3516
rect 564492 3476 564498 3488
rect 565722 3476 565728 3488
rect 565780 3476 565786 3528
rect 568022 3476 568028 3528
rect 568080 3516 568086 3528
rect 569218 3516 569224 3528
rect 568080 3488 569224 3516
rect 568080 3476 568086 3488
rect 569218 3476 569224 3488
rect 569276 3476 569282 3528
rect 571518 3476 571524 3528
rect 571576 3516 571582 3528
rect 572622 3516 572628 3528
rect 571576 3488 572628 3516
rect 571576 3476 571582 3488
rect 572622 3476 572628 3488
rect 572680 3476 572686 3528
rect 573910 3476 573916 3528
rect 573968 3516 573974 3528
rect 575566 3516 575572 3528
rect 573968 3488 575572 3516
rect 573968 3476 573974 3488
rect 575566 3476 575572 3488
rect 575624 3476 575630 3528
rect 576302 3476 576308 3528
rect 576360 3516 576366 3528
rect 576762 3516 576768 3528
rect 576360 3488 576768 3516
rect 576360 3476 576366 3488
rect 576762 3476 576768 3488
rect 576820 3476 576826 3528
rect 577406 3476 577412 3528
rect 577464 3516 577470 3528
rect 578418 3516 578424 3528
rect 577464 3488 578424 3516
rect 577464 3476 577470 3488
rect 578418 3476 578424 3488
rect 578476 3476 578482 3528
rect 483032 3420 489316 3448
rect 489365 3451 489423 3457
rect 489365 3417 489377 3451
rect 489411 3448 489423 3451
rect 512086 3448 512092 3460
rect 489411 3420 512092 3448
rect 489411 3417 489423 3420
rect 489365 3411 489423 3417
rect 512086 3408 512092 3420
rect 512144 3408 512150 3460
rect 514754 3408 514760 3460
rect 514812 3448 514818 3460
rect 530578 3448 530584 3460
rect 514812 3420 530584 3448
rect 514812 3408 514818 3420
rect 530578 3408 530584 3420
rect 530636 3408 530642 3460
rect 554958 3408 554964 3460
rect 555016 3448 555022 3460
rect 556798 3448 556804 3460
rect 555016 3420 556804 3448
rect 555016 3408 555022 3420
rect 556798 3408 556804 3420
rect 556856 3408 556862 3460
rect 559742 3408 559748 3460
rect 559800 3448 559806 3460
rect 560938 3448 560944 3460
rect 559800 3420 560944 3448
rect 559800 3408 559806 3420
rect 560938 3408 560944 3420
rect 560996 3408 561002 3460
rect 570322 3408 570328 3460
rect 570380 3448 570386 3460
rect 574186 3448 574192 3460
rect 570380 3420 574192 3448
rect 570380 3408 570386 3420
rect 574186 3408 574192 3420
rect 574244 3408 574250 3460
rect 471011 3352 474872 3380
rect 471011 3349 471023 3352
rect 470965 3343 471023 3349
rect 478138 3340 478144 3392
rect 478196 3380 478202 3392
rect 501598 3380 501604 3392
rect 478196 3352 501604 3380
rect 478196 3340 478202 3352
rect 501598 3340 501604 3352
rect 501656 3340 501662 3392
rect 502889 3383 502947 3389
rect 502889 3349 502901 3383
rect 502935 3380 502947 3383
rect 508498 3380 508504 3392
rect 502935 3352 508504 3380
rect 502935 3349 502947 3352
rect 502889 3343 502947 3349
rect 508498 3340 508504 3352
rect 508556 3340 508562 3392
rect 530118 3340 530124 3392
rect 530176 3380 530182 3392
rect 531222 3380 531228 3392
rect 530176 3352 531228 3380
rect 530176 3340 530182 3352
rect 531222 3340 531228 3352
rect 531280 3340 531286 3392
rect 536098 3340 536104 3392
rect 536156 3380 536162 3392
rect 540238 3380 540244 3392
rect 536156 3352 540244 3380
rect 536156 3340 536162 3352
rect 540238 3340 540244 3352
rect 540296 3340 540302 3392
rect 553762 3340 553768 3392
rect 553820 3380 553826 3392
rect 561858 3380 561864 3392
rect 553820 3352 561864 3380
rect 553820 3340 553826 3352
rect 561858 3340 561864 3352
rect 561916 3340 561922 3392
rect 466270 3272 466276 3324
rect 466328 3312 466334 3324
rect 468478 3312 468484 3324
rect 466328 3284 468484 3312
rect 466328 3272 466334 3284
rect 468478 3272 468484 3284
rect 468536 3272 468542 3324
rect 476942 3272 476948 3324
rect 477000 3312 477006 3324
rect 497458 3312 497464 3324
rect 477000 3284 497464 3312
rect 477000 3272 477006 3284
rect 497458 3272 497464 3284
rect 497516 3272 497522 3324
rect 529014 3272 529020 3324
rect 529072 3312 529078 3324
rect 537478 3312 537484 3324
rect 529072 3284 537484 3312
rect 529072 3272 529078 3284
rect 537478 3272 537484 3284
rect 537536 3272 537542 3324
rect 562042 3272 562048 3324
rect 562100 3312 562106 3324
rect 566458 3312 566464 3324
rect 562100 3284 566464 3312
rect 562100 3272 562106 3284
rect 566458 3272 566464 3284
rect 566516 3272 566522 3324
rect 469306 3244 469312 3256
rect 462700 3216 469312 3244
rect 462593 3207 462651 3213
rect 469306 3204 469312 3216
rect 469364 3204 469370 3256
rect 474550 3204 474556 3256
rect 474608 3244 474614 3256
rect 480441 3247 480499 3253
rect 480441 3244 480453 3247
rect 474608 3216 480453 3244
rect 474608 3204 474614 3216
rect 480441 3213 480453 3216
rect 480487 3213 480499 3247
rect 480441 3207 480499 3213
rect 480530 3204 480536 3256
rect 480588 3244 480594 3256
rect 489365 3247 489423 3253
rect 489365 3244 489377 3247
rect 480588 3216 489377 3244
rect 480588 3204 480594 3216
rect 489365 3213 489377 3216
rect 489411 3213 489423 3247
rect 489365 3207 489423 3213
rect 569126 3204 569132 3256
rect 569184 3244 569190 3256
rect 572898 3244 572904 3256
rect 569184 3216 572904 3244
rect 569184 3204 569190 3216
rect 572898 3204 572904 3216
rect 572956 3204 572962 3256
rect 338758 3176 338764 3188
rect 302016 3080 305960 3108
rect 306346 3148 338764 3176
rect 302016 3068 302022 3080
rect 306346 3040 306374 3148
rect 338758 3136 338764 3148
rect 338816 3136 338822 3188
rect 340966 3136 340972 3188
rect 341024 3176 341030 3188
rect 416774 3176 416780 3188
rect 341024 3148 416780 3176
rect 341024 3136 341030 3148
rect 416774 3136 416780 3148
rect 416832 3136 416838 3188
rect 422297 3179 422355 3185
rect 422297 3145 422309 3179
rect 422343 3176 422355 3179
rect 426434 3176 426440 3188
rect 422343 3148 426440 3176
rect 422343 3145 422355 3148
rect 422297 3139 422355 3145
rect 426434 3136 426440 3148
rect 426492 3136 426498 3188
rect 428458 3136 428464 3188
rect 428516 3176 428522 3188
rect 472618 3176 472624 3188
rect 428516 3148 472624 3176
rect 428516 3136 428522 3148
rect 472618 3136 472624 3148
rect 472676 3136 472682 3188
rect 473446 3136 473452 3188
rect 473504 3176 473510 3188
rect 482278 3176 482284 3188
rect 473504 3148 482284 3176
rect 473504 3136 473510 3148
rect 482278 3136 482284 3148
rect 482336 3136 482342 3188
rect 532510 3136 532516 3188
rect 532568 3176 532574 3188
rect 538858 3176 538864 3188
rect 532568 3148 538864 3176
rect 532568 3136 532574 3148
rect 538858 3136 538864 3148
rect 538916 3136 538922 3188
rect 539594 3136 539600 3188
rect 539652 3176 539658 3188
rect 543090 3176 543096 3188
rect 539652 3148 543096 3176
rect 539652 3136 539658 3148
rect 543090 3136 543096 3148
rect 543148 3136 543154 3188
rect 552658 3136 552664 3188
rect 552716 3176 552722 3188
rect 555418 3176 555424 3188
rect 552716 3148 555424 3176
rect 552716 3136 552722 3148
rect 555418 3136 555424 3148
rect 555476 3136 555482 3188
rect 563238 3136 563244 3188
rect 563296 3176 563302 3188
rect 565078 3176 565084 3188
rect 563296 3148 565084 3176
rect 563296 3136 563302 3148
rect 565078 3136 565084 3148
rect 565136 3136 565142 3188
rect 583113 3179 583171 3185
rect 583113 3145 583125 3179
rect 583159 3176 583171 3179
rect 583386 3176 583392 3188
rect 583159 3148 583392 3176
rect 583159 3145 583171 3148
rect 583113 3139 583171 3145
rect 583386 3136 583392 3148
rect 583444 3136 583450 3188
rect 307938 3068 307944 3120
rect 307996 3108 308002 3120
rect 311618 3108 311624 3120
rect 307996 3080 311624 3108
rect 307996 3068 308002 3080
rect 311618 3068 311624 3080
rect 311676 3068 311682 3120
rect 316129 3111 316187 3117
rect 316129 3077 316141 3111
rect 316175 3108 316187 3111
rect 324958 3108 324964 3120
rect 316175 3080 324964 3108
rect 316175 3077 316187 3080
rect 316129 3071 316187 3077
rect 324958 3068 324964 3080
rect 325016 3068 325022 3120
rect 325602 3068 325608 3120
rect 325660 3108 325666 3120
rect 370498 3108 370504 3120
rect 325660 3080 370504 3108
rect 325660 3068 325666 3080
rect 370498 3068 370504 3080
rect 370556 3068 370562 3120
rect 376478 3068 376484 3120
rect 376536 3108 376542 3120
rect 382277 3111 382335 3117
rect 382277 3108 382289 3111
rect 376536 3080 382289 3108
rect 376536 3068 376542 3080
rect 382277 3077 382289 3080
rect 382323 3077 382335 3111
rect 382277 3071 382335 3077
rect 394234 3068 394240 3120
rect 394292 3108 394298 3120
rect 396718 3108 396724 3120
rect 394292 3080 396724 3108
rect 394292 3068 394298 3080
rect 396718 3068 396724 3080
rect 396776 3068 396782 3120
rect 404541 3111 404599 3117
rect 404541 3077 404553 3111
rect 404587 3108 404599 3111
rect 411254 3108 411260 3120
rect 404587 3080 411260 3108
rect 404587 3077 404599 3080
rect 404541 3071 404599 3077
rect 411254 3068 411260 3080
rect 411312 3068 411318 3120
rect 411898 3068 411904 3120
rect 411956 3108 411962 3120
rect 460198 3108 460204 3120
rect 411956 3080 460204 3108
rect 411956 3068 411962 3080
rect 460198 3068 460204 3080
rect 460256 3068 460262 3120
rect 463970 3068 463976 3120
rect 464028 3108 464034 3120
rect 483658 3108 483664 3120
rect 464028 3080 483664 3108
rect 464028 3068 464034 3080
rect 483658 3068 483664 3080
rect 483716 3068 483722 3120
rect 301516 3012 306374 3040
rect 318518 3000 318524 3052
rect 318576 3040 318582 3052
rect 360838 3040 360844 3052
rect 318576 3012 360844 3040
rect 318576 3000 318582 3012
rect 360838 3000 360844 3012
rect 360896 3000 360902 3052
rect 387150 3000 387156 3052
rect 387208 3040 387214 3052
rect 387702 3040 387708 3052
rect 387208 3012 387708 3040
rect 387208 3000 387214 3012
rect 387702 3000 387708 3012
rect 387760 3000 387766 3052
rect 396534 3000 396540 3052
rect 396592 3040 396598 3052
rect 402333 3043 402391 3049
rect 402333 3040 402345 3043
rect 396592 3012 402345 3040
rect 396592 3000 396598 3012
rect 402333 3009 402345 3012
rect 402379 3009 402391 3043
rect 402333 3003 402391 3009
rect 409598 3000 409604 3052
rect 409656 3040 409662 3052
rect 413278 3040 413284 3052
rect 409656 3012 413284 3040
rect 409656 3000 409662 3012
rect 413278 3000 413284 3012
rect 413336 3000 413342 3052
rect 417878 3000 417884 3052
rect 417936 3040 417942 3052
rect 422941 3043 422999 3049
rect 422941 3040 422953 3043
rect 417936 3012 422953 3040
rect 417936 3000 417942 3012
rect 422941 3009 422953 3012
rect 422987 3009 422999 3043
rect 422941 3003 422999 3009
rect 439130 3000 439136 3052
rect 439188 3040 439194 3052
rect 474090 3040 474096 3052
rect 439188 3012 474096 3040
rect 439188 3000 439194 3012
rect 474090 3000 474096 3012
rect 474148 3000 474154 3052
rect 486418 3000 486424 3052
rect 486476 3040 486482 3052
rect 487062 3040 487068 3052
rect 486476 3012 487068 3040
rect 486476 3000 486482 3012
rect 487062 3000 487068 3012
rect 487120 3000 487126 3052
rect 494698 3000 494704 3052
rect 494756 3040 494762 3052
rect 495342 3040 495348 3052
rect 494756 3012 495348 3040
rect 494756 3000 494762 3012
rect 495342 3000 495348 3012
rect 495400 3000 495406 3052
rect 578602 3000 578608 3052
rect 578660 3040 578666 3052
rect 579614 3040 579620 3052
rect 578660 3012 579620 3040
rect 578660 3000 578666 3012
rect 579614 3000 579620 3012
rect 579672 3000 579678 3052
rect 110564 2944 113174 2972
rect 110564 2932 110570 2944
rect 114002 2932 114008 2984
rect 114060 2972 114066 2984
rect 114462 2972 114468 2984
rect 114060 2944 114468 2972
rect 114060 2932 114066 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 116394 2932 116400 2984
rect 116452 2972 116458 2984
rect 117222 2972 117228 2984
rect 116452 2944 117228 2972
rect 116452 2932 116458 2944
rect 117222 2932 117228 2944
rect 117280 2932 117286 2984
rect 118786 2932 118792 2984
rect 118844 2972 118850 2984
rect 119798 2972 119804 2984
rect 118844 2944 119804 2972
rect 118844 2932 118850 2944
rect 119798 2932 119804 2944
rect 119856 2932 119862 2984
rect 122282 2932 122288 2984
rect 122340 2972 122346 2984
rect 122742 2972 122748 2984
rect 122340 2944 122748 2972
rect 122340 2932 122346 2944
rect 122742 2932 122748 2944
rect 122800 2932 122806 2984
rect 123478 2932 123484 2984
rect 123536 2972 123542 2984
rect 124122 2972 124128 2984
rect 123536 2944 124128 2972
rect 123536 2932 123542 2944
rect 124122 2932 124128 2944
rect 124180 2932 124186 2984
rect 125870 2932 125876 2984
rect 125928 2972 125934 2984
rect 126882 2972 126888 2984
rect 125928 2944 126888 2972
rect 125928 2932 125934 2944
rect 126882 2932 126888 2944
rect 126940 2932 126946 2984
rect 232498 2972 232504 2984
rect 127636 2944 232504 2972
rect 105538 2904 105544 2916
rect 93826 2876 105544 2904
rect 105538 2864 105544 2876
rect 105596 2864 105602 2916
rect 117590 2864 117596 2916
rect 117648 2904 117654 2916
rect 127636 2904 127664 2944
rect 232498 2932 232504 2944
rect 232556 2932 232562 2984
rect 309042 2932 309048 2984
rect 309100 2972 309106 2984
rect 329098 2972 329104 2984
rect 309100 2944 329104 2972
rect 309100 2932 309106 2944
rect 329098 2932 329104 2944
rect 329156 2932 329162 2984
rect 332686 2932 332692 2984
rect 332744 2972 332750 2984
rect 356698 2972 356704 2984
rect 332744 2944 356704 2972
rect 332744 2932 332750 2944
rect 356698 2932 356704 2944
rect 356756 2932 356762 2984
rect 357526 2932 357532 2984
rect 357584 2972 357590 2984
rect 359458 2972 359464 2984
rect 357584 2944 359464 2972
rect 357584 2932 357590 2944
rect 359458 2932 359464 2944
rect 359516 2932 359522 2984
rect 364610 2932 364616 2984
rect 364668 2972 364674 2984
rect 376018 2972 376024 2984
rect 364668 2944 376024 2972
rect 364668 2932 364674 2944
rect 376018 2932 376024 2944
rect 376076 2932 376082 2984
rect 413005 2975 413063 2981
rect 413005 2941 413017 2975
rect 413051 2972 413063 2975
rect 420914 2972 420920 2984
rect 413051 2944 420920 2972
rect 413051 2941 413063 2944
rect 413005 2935 413063 2941
rect 420914 2932 420920 2944
rect 420972 2932 420978 2984
rect 431957 2975 432015 2981
rect 431957 2941 431969 2975
rect 432003 2972 432015 2975
rect 442258 2972 442264 2984
rect 432003 2944 442264 2972
rect 432003 2941 432015 2944
rect 431957 2935 432015 2941
rect 442258 2932 442264 2944
rect 442316 2932 442322 2984
rect 442626 2932 442632 2984
rect 442684 2972 442690 2984
rect 476758 2972 476764 2984
rect 442684 2944 476764 2972
rect 442684 2932 442690 2944
rect 476758 2932 476764 2944
rect 476816 2932 476822 2984
rect 557350 2932 557356 2984
rect 557408 2972 557414 2984
rect 558178 2972 558184 2984
rect 557408 2944 558184 2972
rect 557408 2932 557414 2944
rect 558178 2932 558184 2944
rect 558236 2932 558242 2984
rect 233878 2904 233884 2916
rect 117648 2876 127664 2904
rect 128096 2876 233884 2904
rect 117648 2864 117654 2876
rect 124674 2796 124680 2848
rect 124732 2836 124738 2848
rect 128096 2836 128124 2876
rect 233878 2864 233884 2876
rect 233936 2864 233942 2916
rect 315022 2864 315028 2916
rect 315080 2904 315086 2916
rect 318058 2904 318064 2916
rect 315080 2876 318064 2904
rect 315080 2864 315086 2876
rect 318058 2864 318064 2876
rect 318116 2864 318122 2916
rect 329190 2864 329196 2916
rect 329248 2904 329254 2916
rect 340049 2907 340107 2913
rect 329248 2876 340000 2904
rect 329248 2864 329254 2876
rect 124732 2808 128124 2836
rect 124732 2796 124738 2808
rect 131758 2796 131764 2848
rect 131816 2836 131822 2848
rect 132402 2836 132408 2848
rect 131816 2808 132408 2836
rect 131816 2796 131822 2808
rect 132402 2796 132408 2808
rect 132460 2796 132466 2848
rect 132954 2796 132960 2848
rect 133012 2836 133018 2848
rect 133782 2836 133788 2848
rect 133012 2808 133788 2836
rect 133012 2796 133018 2808
rect 133782 2796 133788 2808
rect 133840 2796 133846 2848
rect 134150 2796 134156 2848
rect 134208 2836 134214 2848
rect 135162 2836 135168 2848
rect 134208 2808 135168 2836
rect 134208 2796 134214 2808
rect 135162 2796 135168 2808
rect 135220 2796 135226 2848
rect 140038 2796 140044 2848
rect 140096 2836 140102 2848
rect 140682 2836 140688 2848
rect 140096 2808 140688 2836
rect 140096 2796 140102 2808
rect 140682 2796 140688 2808
rect 140740 2796 140746 2848
rect 141234 2796 141240 2848
rect 141292 2836 141298 2848
rect 142062 2836 142068 2848
rect 141292 2808 142068 2836
rect 141292 2796 141298 2808
rect 142062 2796 142068 2808
rect 142120 2796 142126 2848
rect 143534 2796 143540 2848
rect 143592 2836 143598 2848
rect 144822 2836 144828 2848
rect 143592 2808 144828 2836
rect 143592 2796 143598 2808
rect 144822 2796 144828 2808
rect 144880 2796 144886 2848
rect 147122 2796 147128 2848
rect 147180 2836 147186 2848
rect 147582 2836 147588 2848
rect 147180 2808 147588 2836
rect 147180 2796 147186 2808
rect 147582 2796 147588 2808
rect 147640 2796 147646 2848
rect 148318 2796 148324 2848
rect 148376 2836 148382 2848
rect 148962 2836 148968 2848
rect 148376 2808 148968 2836
rect 148376 2796 148382 2808
rect 148962 2796 148968 2808
rect 149020 2796 149026 2848
rect 150618 2796 150624 2848
rect 150676 2836 150682 2848
rect 151722 2836 151728 2848
rect 150676 2808 151728 2836
rect 150676 2796 150682 2808
rect 151722 2796 151728 2808
rect 151780 2796 151786 2848
rect 151814 2796 151820 2848
rect 151872 2836 151878 2848
rect 153102 2836 153108 2848
rect 151872 2808 153108 2836
rect 151872 2796 151878 2808
rect 153102 2796 153108 2808
rect 153160 2796 153166 2848
rect 155402 2796 155408 2848
rect 155460 2836 155466 2848
rect 155862 2836 155868 2848
rect 155460 2808 155868 2836
rect 155460 2796 155466 2808
rect 155862 2796 155868 2808
rect 155920 2796 155926 2848
rect 157794 2796 157800 2848
rect 157852 2836 157858 2848
rect 158622 2836 158628 2848
rect 157852 2808 158628 2836
rect 157852 2796 157858 2808
rect 158622 2796 158628 2808
rect 158680 2796 158686 2848
rect 164878 2796 164884 2848
rect 164936 2836 164942 2848
rect 165522 2836 165528 2848
rect 164936 2808 165528 2836
rect 164936 2796 164942 2808
rect 165522 2796 165528 2808
rect 165580 2796 165586 2848
rect 168374 2796 168380 2848
rect 168432 2836 168438 2848
rect 169662 2836 169668 2848
rect 168432 2808 169668 2836
rect 168432 2796 168438 2808
rect 169662 2796 169668 2808
rect 169720 2796 169726 2848
rect 171962 2796 171968 2848
rect 172020 2836 172026 2848
rect 172422 2836 172428 2848
rect 172020 2808 172428 2836
rect 172020 2796 172026 2808
rect 172422 2796 172428 2808
rect 172480 2796 172486 2848
rect 175458 2796 175464 2848
rect 175516 2836 175522 2848
rect 176562 2836 176568 2848
rect 175516 2808 176568 2836
rect 175516 2796 175522 2808
rect 176562 2796 176568 2808
rect 176620 2796 176626 2848
rect 181349 2839 181407 2845
rect 181349 2805 181361 2839
rect 181395 2836 181407 2839
rect 189166 2836 189172 2848
rect 181395 2808 189172 2836
rect 181395 2805 181407 2808
rect 181349 2799 181407 2805
rect 189166 2796 189172 2808
rect 189224 2796 189230 2848
rect 229830 2796 229836 2848
rect 229888 2836 229894 2848
rect 231394 2836 231400 2848
rect 229888 2808 231400 2836
rect 229888 2796 229894 2808
rect 231394 2796 231400 2808
rect 231452 2796 231458 2848
rect 325697 2839 325755 2845
rect 325697 2805 325709 2839
rect 325743 2836 325755 2839
rect 332045 2839 332103 2845
rect 332045 2836 332057 2839
rect 325743 2808 332057 2836
rect 325743 2805 325755 2808
rect 325697 2799 325755 2805
rect 332045 2805 332057 2808
rect 332091 2805 332103 2839
rect 332045 2799 332103 2805
rect 333882 2796 333888 2848
rect 333940 2836 333946 2848
rect 339865 2839 339923 2845
rect 339865 2836 339877 2839
rect 333940 2808 339877 2836
rect 333940 2796 333946 2808
rect 339865 2805 339877 2808
rect 339911 2805 339923 2839
rect 339865 2799 339923 2805
rect 339972 2768 340000 2876
rect 340049 2873 340061 2907
rect 340095 2904 340107 2907
rect 347038 2904 347044 2916
rect 340095 2876 347044 2904
rect 340095 2873 340107 2876
rect 340049 2867 340107 2873
rect 347038 2864 347044 2876
rect 347096 2864 347102 2916
rect 388254 2864 388260 2916
rect 388312 2904 388318 2916
rect 389818 2904 389824 2916
rect 388312 2876 389824 2904
rect 388312 2864 388318 2876
rect 389818 2864 389824 2876
rect 389876 2864 389882 2916
rect 444929 2907 444987 2913
rect 444929 2873 444941 2907
rect 444975 2904 444987 2907
rect 453206 2904 453212 2916
rect 444975 2876 453212 2904
rect 444975 2873 444987 2876
rect 444929 2867 444987 2873
rect 453206 2864 453212 2876
rect 453264 2864 453270 2916
rect 453298 2864 453304 2916
rect 453356 2904 453362 2916
rect 475378 2904 475384 2916
rect 453356 2876 475384 2904
rect 453356 2864 453362 2876
rect 475378 2864 475384 2876
rect 475436 2864 475442 2916
rect 572714 2864 572720 2916
rect 572772 2904 572778 2916
rect 574002 2904 574008 2916
rect 572772 2876 574008 2904
rect 572772 2864 572778 2876
rect 574002 2864 574008 2876
rect 574060 2864 574066 2916
rect 341518 2836 341524 2848
rect 340248 2808 341524 2836
rect 340248 2768 340276 2808
rect 341518 2796 341524 2808
rect 341576 2796 341582 2848
rect 434438 2796 434444 2848
rect 434496 2836 434502 2848
rect 447870 2836 447876 2848
rect 434496 2808 447876 2836
rect 434496 2796 434502 2808
rect 447870 2796 447876 2808
rect 447928 2796 447934 2848
rect 448606 2796 448612 2848
rect 448664 2836 448670 2848
rect 461486 2836 461492 2848
rect 448664 2808 461492 2836
rect 448664 2796 448670 2808
rect 461486 2796 461492 2808
rect 461544 2796 461550 2848
rect 339972 2740 340276 2768
<< via1 >>
rect 15844 703740 15896 703792
rect 552940 703740 552992 703792
rect 22744 703672 22796 703724
rect 563520 703672 563572 703724
rect 363512 703604 363564 703656
rect 429660 703604 429712 703656
rect 300308 703536 300360 703588
rect 384580 703536 384632 703588
rect 374552 703468 374604 703520
rect 577044 703468 577096 703520
rect 182180 703400 182232 703452
rect 437204 703400 437256 703452
rect 349436 703332 349488 703384
rect 543464 703332 543516 703384
rect 182272 703264 182324 703316
rect 447692 703264 447744 703316
rect 182364 703196 182416 703248
rect 458180 703196 458232 703248
rect 182456 703128 182508 703180
rect 468760 703128 468812 703180
rect 182548 703060 182600 703112
rect 479248 703060 479300 703112
rect 182640 702992 182692 703044
rect 489828 702992 489880 703044
rect 182732 702924 182784 702976
rect 500316 702924 500368 702976
rect 258172 702856 258224 702908
rect 254676 702788 254728 702840
rect 226616 702720 226668 702772
rect 180064 702652 180116 702704
rect 542452 702652 542504 702704
rect 219624 702584 219676 702636
rect 300308 702516 300360 702568
rect 375380 702516 375432 702568
rect 404360 702516 404412 702568
rect 409052 702516 409104 702568
rect 365720 702448 365772 702500
rect 369676 702491 369728 702500
rect 369676 702457 369685 702491
rect 369685 702457 369719 702491
rect 369719 702457 369728 702491
rect 369676 702448 369728 702457
rect 370504 702448 370556 702500
rect 413652 702448 413704 702500
rect 35164 702380 35216 702432
rect 486332 702380 486384 702432
rect 18604 702312 18656 702364
rect 475752 702312 475804 702364
rect 14464 702244 14516 702296
rect 472256 702244 472308 702296
rect 289820 702176 289872 702228
rect 333980 702176 334032 702228
rect 338948 702176 339000 702228
rect 427636 702176 427688 702228
rect 314384 702108 314436 702160
rect 418068 702108 418120 702160
rect 268752 702040 268804 702092
rect 374552 702040 374604 702092
rect 374644 702040 374696 702092
rect 556436 702040 556488 702092
rect 328368 701972 328420 702024
rect 583760 701972 583812 702024
rect 324872 701904 324924 701956
rect 583852 701904 583904 701956
rect 307300 701836 307352 701888
rect 583576 701836 583628 701888
rect 304080 701768 304132 701820
rect 582564 701768 582616 701820
rect 181812 701700 181864 701752
rect 182088 701632 182140 701684
rect 297088 701700 297140 701752
rect 583392 701700 583444 701752
rect 181904 701564 181956 701616
rect 201684 701632 201736 701684
rect 293592 701632 293644 701684
rect 583484 701632 583536 701684
rect 191196 701564 191248 701616
rect 286600 701564 286652 701616
rect 583208 701564 583260 701616
rect 183008 701496 183060 701548
rect 205180 701496 205232 701548
rect 282828 701496 282880 701548
rect 583300 701496 583352 701548
rect 182916 701428 182968 701480
rect 208676 701428 208728 701480
rect 279608 701428 279660 701480
rect 583116 701428 583168 701480
rect 137284 701360 137336 701412
rect 244004 701360 244056 701412
rect 275928 701360 275980 701412
rect 582932 701360 582984 701412
rect 39304 701292 39356 701344
rect 247868 701292 247920 701344
rect 272616 701292 272668 701344
rect 583024 701292 583076 701344
rect 32404 701224 32456 701276
rect 482468 701224 482520 701276
rect 183100 701156 183152 701208
rect 194692 701156 194744 701208
rect 362224 701199 362276 701208
rect 362224 701165 362233 701199
rect 362233 701165 362267 701199
rect 362267 701165 362276 701199
rect 362224 701156 362276 701165
rect 362960 701156 363012 701208
rect 364984 701199 365036 701208
rect 364984 701165 364993 701199
rect 364993 701165 365027 701199
rect 365027 701165 365036 701199
rect 364984 701156 365036 701165
rect 367100 701156 367152 701208
rect 391112 701199 391164 701208
rect 391112 701165 391121 701199
rect 391121 701165 391155 701199
rect 391155 701165 391164 701199
rect 391112 701156 391164 701165
rect 532240 701156 532292 701208
rect 535552 701156 535604 701208
rect 181996 701088 182048 701140
rect 187700 701088 187752 701140
rect 198188 701088 198240 701140
rect 316132 701131 316184 701140
rect 316132 701097 316141 701131
rect 316141 701097 316175 701131
rect 316175 701097 316184 701131
rect 316132 701088 316184 701097
rect 182824 701020 182876 701072
rect 184204 701020 184256 701072
rect 202788 701063 202840 701072
rect 202788 701029 202797 701063
rect 202797 701029 202831 701063
rect 202831 701029 202840 701063
rect 202788 701020 202840 701029
rect 262036 701063 262088 701072
rect 262036 701029 262045 701063
rect 262045 701029 262079 701063
rect 262079 701029 262088 701063
rect 262036 701020 262088 701029
rect 265624 701063 265676 701072
rect 265624 701029 265633 701063
rect 265633 701029 265667 701063
rect 265667 701029 265676 701063
rect 265624 701020 265676 701029
rect 267648 701063 267700 701072
rect 267648 701029 267657 701063
rect 267657 701029 267691 701063
rect 267691 701029 267700 701063
rect 267648 701020 267700 701029
rect 283840 701063 283892 701072
rect 283840 701029 283849 701063
rect 283849 701029 283883 701063
rect 283883 701029 283892 701063
rect 283840 701020 283892 701029
rect 318248 701063 318300 701072
rect 318248 701029 318257 701063
rect 318257 701029 318291 701063
rect 318291 701029 318300 701063
rect 318248 701020 318300 701029
rect 137836 700952 137888 701004
rect 332508 701020 332560 701072
rect 335728 701088 335780 701140
rect 365812 701088 365864 701140
rect 369492 701088 369544 701140
rect 373816 701131 373868 701140
rect 373816 701097 373825 701131
rect 373825 701097 373859 701131
rect 373859 701097 373868 701131
rect 373816 701088 373868 701097
rect 374092 701131 374144 701140
rect 374092 701097 374101 701131
rect 374101 701097 374135 701131
rect 374135 701097 374144 701131
rect 374092 701088 374144 701097
rect 377220 701131 377272 701140
rect 377220 701097 377229 701131
rect 377229 701097 377263 701131
rect 377263 701097 377272 701131
rect 377220 701088 377272 701097
rect 387800 701131 387852 701140
rect 387800 701097 387809 701131
rect 387809 701097 387843 701131
rect 387843 701097 387852 701131
rect 387800 701088 387852 701097
rect 391204 701131 391256 701140
rect 391204 701097 391213 701131
rect 391213 701097 391247 701131
rect 391247 701097 391256 701131
rect 391204 701088 391256 701097
rect 397460 701131 397512 701140
rect 397460 701097 397469 701131
rect 397469 701097 397503 701131
rect 397503 701097 397512 701131
rect 397460 701088 397512 701097
rect 333244 701063 333296 701072
rect 333244 701029 333253 701063
rect 333253 701029 333287 701063
rect 333287 701029 333296 701063
rect 333244 701020 333296 701029
rect 349068 701063 349120 701072
rect 349068 701029 349077 701063
rect 349077 701029 349111 701063
rect 349111 701029 349120 701063
rect 349068 701020 349120 701029
rect 356704 701063 356756 701072
rect 356704 701029 356713 701063
rect 356713 701029 356747 701063
rect 356747 701029 356756 701063
rect 356704 701020 356756 701029
rect 360108 701020 360160 701072
rect 398196 701063 398248 701072
rect 398196 701029 398205 701063
rect 398205 701029 398239 701063
rect 398239 701029 398248 701063
rect 398196 701020 398248 701029
rect 401692 701063 401744 701072
rect 401692 701029 401701 701063
rect 401701 701029 401735 701063
rect 401735 701029 401744 701063
rect 401692 701020 401744 701029
rect 404360 701020 404412 701072
rect 419724 701063 419776 701072
rect 419724 701029 419733 701063
rect 419733 701029 419767 701063
rect 419767 701029 419776 701063
rect 419724 701020 419776 701029
rect 422852 701063 422904 701072
rect 422852 701029 422861 701063
rect 422861 701029 422895 701063
rect 422895 701029 422904 701063
rect 422852 701020 422904 701029
rect 429844 701063 429896 701072
rect 429844 701029 429853 701063
rect 429853 701029 429887 701063
rect 429887 701029 429896 701063
rect 429844 701020 429896 701029
rect 433340 701063 433392 701072
rect 433340 701029 433349 701063
rect 433349 701029 433383 701063
rect 433383 701029 433392 701063
rect 433340 701020 433392 701029
rect 440332 701063 440384 701072
rect 440332 701029 440341 701063
rect 440341 701029 440375 701063
rect 440375 701029 440384 701063
rect 440332 701020 440384 701029
rect 443828 701063 443880 701072
rect 443828 701029 443837 701063
rect 443837 701029 443871 701063
rect 443871 701029 443880 701063
rect 443828 701020 443880 701029
rect 450820 701063 450872 701072
rect 450820 701029 450829 701063
rect 450829 701029 450863 701063
rect 450863 701029 450872 701063
rect 450820 701020 450872 701029
rect 454316 701063 454368 701072
rect 454316 701029 454325 701063
rect 454325 701029 454359 701063
rect 454359 701029 454368 701063
rect 454316 701020 454368 701029
rect 461492 701063 461544 701072
rect 461492 701029 461501 701063
rect 461501 701029 461535 701063
rect 461535 701029 461544 701063
rect 461492 701020 461544 701029
rect 462320 701063 462372 701072
rect 462320 701029 462329 701063
rect 462329 701029 462363 701063
rect 462363 701029 462372 701063
rect 462320 701020 462372 701029
rect 465080 701063 465132 701072
rect 465080 701029 465089 701063
rect 465089 701029 465123 701063
rect 465123 701029 465132 701063
rect 465080 701020 465132 701029
rect 478512 701020 478564 701072
rect 566740 701020 566792 701072
rect 577872 701020 577924 701072
rect 61384 700544 61436 700596
rect 36544 700476 36596 700528
rect 583668 700476 583720 700528
rect 582748 700408 582800 700460
rect 582840 700340 582892 700392
rect 89168 700272 89220 700324
rect 72976 700204 73028 700256
rect 24308 700136 24360 700188
rect 32496 700068 32548 700120
rect 35256 700000 35308 700052
rect 8116 699932 8168 699984
rect 40776 699864 40828 699916
rect 18696 699796 18748 699848
rect 14556 699728 14608 699780
rect 33876 699660 33928 699712
rect 3516 684428 3568 684480
rect 182180 684428 182232 684480
rect 3056 671984 3108 672036
rect 18696 671984 18748 672036
rect 3516 658180 3568 658232
rect 14556 658180 14608 658232
rect 3240 633360 3292 633412
rect 182272 633360 182324 633412
rect 3332 619556 3384 619608
rect 35256 619556 35308 619608
rect 3240 607112 3292 607164
rect 32496 607112 32548 607164
rect 3148 580932 3200 580984
rect 182364 580932 182416 580984
rect 3516 567128 3568 567180
rect 40776 567128 40828 567180
rect 3516 554684 3568 554736
rect 33876 554684 33928 554736
rect 2872 528504 2924 528556
rect 182456 528504 182508 528556
rect 3516 516060 3568 516112
rect 18604 516060 18656 516112
rect 3516 502256 3568 502308
rect 14464 502256 14516 502308
rect 3516 476008 3568 476060
rect 182548 476008 182600 476060
rect 3240 463632 3292 463684
rect 35164 463632 35216 463684
rect 3332 449828 3384 449880
rect 32404 449828 32456 449880
rect 3516 423580 3568 423632
rect 182640 423580 182692 423632
rect 2964 411204 3016 411256
rect 25504 411204 25556 411256
rect 3240 398760 3292 398812
rect 17224 398760 17276 398812
rect 3516 372512 3568 372564
rect 182732 372512 182784 372564
rect 3332 358708 3384 358760
rect 29644 358708 29696 358760
rect 3148 346332 3200 346384
rect 177304 346332 177356 346384
rect 3332 318792 3384 318844
rect 182732 318792 182784 318844
rect 3516 306280 3568 306332
rect 33784 306280 33836 306332
rect 182824 302948 182876 303000
rect 181812 302880 181864 302932
rect 580264 302404 580316 302456
rect 580356 302336 580408 302388
rect 182180 299480 182232 299532
rect 183192 299480 183244 299532
rect 183560 299480 183612 299532
rect 184388 299480 184440 299532
rect 351920 299480 351972 299532
rect 352380 299480 352432 299532
rect 353392 299480 353444 299532
rect 354036 299480 354088 299532
rect 367100 299480 367152 299532
rect 367836 299480 367888 299532
rect 440240 299480 440292 299532
rect 440884 299480 440936 299532
rect 107568 299412 107620 299464
rect 256148 299412 256200 299464
rect 258080 299412 258132 299464
rect 265072 299412 265124 299464
rect 293500 299412 293552 299464
rect 296076 299412 296128 299464
rect 313004 299412 313056 299464
rect 335360 299412 335412 299464
rect 336188 299412 336240 299464
rect 338120 299412 338172 299464
rect 338580 299412 338632 299464
rect 339500 299412 339552 299464
rect 340236 299412 340288 299464
rect 414388 299412 414440 299464
rect 416688 299412 416740 299464
rect 103428 299344 103480 299396
rect 253756 299344 253808 299396
rect 90364 299276 90416 299328
rect 244004 299276 244056 299328
rect 246948 299276 247000 299328
rect 248052 299276 248104 299328
rect 253296 299276 253348 299328
rect 273168 299344 273220 299396
rect 274088 299344 274140 299396
rect 317880 299344 317932 299396
rect 331864 299344 331916 299396
rect 409512 299344 409564 299396
rect 410524 299344 410576 299396
rect 416044 299344 416096 299396
rect 420920 299344 420972 299396
rect 421380 299344 421432 299396
rect 467104 299412 467156 299464
rect 474004 299412 474056 299464
rect 479340 299412 479392 299464
rect 493876 299412 493928 299464
rect 501236 299412 501288 299464
rect 523132 299412 523184 299464
rect 526444 299412 526496 299464
rect 541808 299412 541860 299464
rect 547144 299412 547196 299464
rect 557172 299412 557224 299464
rect 467932 299344 467984 299396
rect 298376 299276 298428 299328
rect 300124 299276 300176 299328
rect 308128 299276 308180 299328
rect 313280 299276 313332 299328
rect 314292 299276 314344 299328
rect 320180 299276 320232 299328
rect 320732 299276 320784 299328
rect 325700 299276 325752 299328
rect 326436 299276 326488 299328
rect 327724 299276 327776 299328
rect 404636 299276 404688 299328
rect 408408 299276 408460 299328
rect 463056 299276 463108 299328
rect 467748 299276 467800 299328
rect 469220 299276 469272 299328
rect 470140 299276 470192 299328
rect 472624 299344 472676 299396
rect 476856 299344 476908 299396
rect 478144 299344 478196 299396
rect 506112 299344 506164 299396
rect 507768 299344 507820 299396
rect 530400 299344 530452 299396
rect 530584 299344 530636 299396
rect 536104 299344 536156 299396
rect 503628 299276 503680 299328
rect 504364 299276 504416 299328
rect 506848 299276 506900 299328
rect 522396 299276 522448 299328
rect 524696 299276 524748 299328
rect 525156 299276 525208 299328
rect 527180 299276 527232 299328
rect 529296 299276 529348 299328
rect 531228 299276 531280 299328
rect 533988 299276 534040 299328
rect 549076 299344 549128 299396
rect 558184 299344 558236 299396
rect 565268 299344 565320 299396
rect 569224 299344 569276 299396
rect 572628 299344 572680 299396
rect 546684 299276 546736 299328
rect 548524 299276 548576 299328
rect 558000 299276 558052 299328
rect 560944 299276 560996 299328
rect 566924 299276 566976 299328
rect 574008 299276 574060 299328
rect 575848 299276 575900 299328
rect 582380 299276 582432 299328
rect 50344 299208 50396 299260
rect 214748 299208 214800 299260
rect 232504 299208 232556 299260
rect 263508 299208 263560 299260
rect 263692 299208 263744 299260
rect 274824 299208 274876 299260
rect 281356 299208 281408 299260
rect 283748 299208 283800 299260
rect 285680 299208 285732 299260
rect 286692 299208 286744 299260
rect 355968 299208 356020 299260
rect 357440 299208 357492 299260
rect 358084 299208 358136 299260
rect 358820 299208 358872 299260
rect 359740 299208 359792 299260
rect 362224 299208 362276 299260
rect 363236 299208 363288 299260
rect 429016 299208 429068 299260
rect 430580 299208 430632 299260
rect 431132 299208 431184 299260
rect 477684 299208 477736 299260
rect 478236 299208 478288 299260
rect 480076 299208 480128 299260
rect 480168 299208 480220 299260
rect 484952 299208 485004 299260
rect 493324 299208 493376 299260
rect 496360 299208 496412 299260
rect 519084 299208 519136 299260
rect 519544 299208 519596 299260
rect 523960 299208 524012 299260
rect 539324 299208 539376 299260
rect 540244 299208 540296 299260
rect 550732 299208 550784 299260
rect 551928 299208 551980 299260
rect 561220 299208 561272 299260
rect 572628 299208 572680 299260
rect 575020 299208 575072 299260
rect 35164 299140 35216 299192
rect 195980 299140 196032 299192
rect 196532 299140 196584 299192
rect 201500 299140 201552 299192
rect 202236 299140 202288 299192
rect 220084 299140 220136 299192
rect 241612 299140 241664 299192
rect 246488 299140 246540 299192
rect 300768 299140 300820 299192
rect 312176 299140 312228 299192
rect 312544 299140 312596 299192
rect 319444 299140 319496 299192
rect 322204 299140 322256 299192
rect 399392 299140 399444 299192
rect 399484 299140 399536 299192
rect 402244 299140 402296 299192
rect 456064 299140 456116 299192
rect 460664 299140 460716 299192
rect 497188 299140 497240 299192
rect 503628 299140 503680 299192
rect 526352 299140 526404 299192
rect 527088 299140 527140 299192
rect 544200 299140 544252 299192
rect 544384 299140 544436 299192
rect 555332 299140 555384 299192
rect 555424 299140 555476 299192
rect 562048 299140 562100 299192
rect 43444 299072 43496 299124
rect 209964 299072 210016 299124
rect 217324 299072 217376 299124
rect 239128 299072 239180 299124
rect 253204 299072 253256 299124
rect 295892 299072 295944 299124
rect 295984 299072 296036 299124
rect 33784 299004 33836 299056
rect 205088 299004 205140 299056
rect 227076 299004 227128 299056
rect 258632 299004 258684 299056
rect 262864 299004 262916 299056
rect 279700 299004 279752 299056
rect 282184 299004 282236 299056
rect 370596 299004 370648 299056
rect 371884 299004 371936 299056
rect 372988 299004 373040 299056
rect 373908 299004 373960 299056
rect 29644 298936 29696 298988
rect 200212 298936 200264 298988
rect 214564 298936 214616 298988
rect 234252 298936 234304 298988
rect 234528 298936 234580 298988
rect 268384 298936 268436 298988
rect 268844 298936 268896 298988
rect 280988 298936 281040 298988
rect 284944 298936 284996 298988
rect 375472 298936 375524 298988
rect 376760 299072 376812 299124
rect 377588 299072 377640 299124
rect 380164 299072 380216 299124
rect 442816 299072 442868 299124
rect 443644 299072 443696 299124
rect 445208 299072 445260 299124
rect 449164 299072 449216 299124
rect 450084 299072 450136 299124
rect 491484 299072 491536 299124
rect 493968 299072 494020 299124
rect 521476 299072 521528 299124
rect 528008 299072 528060 299124
rect 540152 299072 540204 299124
rect 435364 299004 435416 299056
rect 436284 299004 436336 299056
rect 436744 299004 436796 299056
rect 437940 299004 437992 299056
rect 438124 299004 438176 299056
rect 482560 299004 482612 299056
rect 485688 299004 485740 299056
rect 515312 299004 515364 299056
rect 515404 299004 515456 299056
rect 535276 299004 535328 299056
rect 536196 299004 536248 299056
rect 543372 299072 543424 299124
rect 545028 299072 545080 299124
rect 556344 299072 556396 299124
rect 543004 299004 543056 299056
rect 554780 299004 554832 299056
rect 380348 298936 380400 298988
rect 380808 298936 380860 298988
rect 442264 298936 442316 298988
rect 446036 298936 446088 298988
rect 449808 298936 449860 298988
rect 487436 298936 487488 298988
rect 489828 298936 489880 298988
rect 518256 298936 518308 298988
rect 518808 298936 518860 298988
rect 538496 298936 538548 298988
rect 540888 298936 540940 298988
rect 553952 298936 554004 298988
rect 556804 298936 556856 298988
rect 563704 298936 563756 298988
rect 18604 298868 18656 298920
rect 192852 298868 192904 298920
rect 199384 298868 199436 298920
rect 211804 298868 211856 298920
rect 224500 298868 224552 298920
rect 17224 298800 17276 298852
rect 193680 298800 193732 298852
rect 210424 298800 210476 298852
rect 219624 298800 219676 298852
rect 224224 298800 224276 298852
rect 251272 298868 251324 298920
rect 255964 298868 256016 298920
rect 246396 298800 246448 298852
rect 249064 298800 249116 298852
rect 346216 298800 346268 298852
rect 347044 298868 347096 298920
rect 348700 298868 348752 298920
rect 351828 298868 351880 298920
rect 424140 298868 424192 298920
rect 430488 298868 430540 298920
rect 351092 298800 351144 298852
rect 419264 298800 419316 298852
rect 424968 298800 425020 298852
rect 474464 298868 474516 298920
rect 476764 298868 476816 298920
rect 486608 298868 486660 298920
rect 487068 298868 487120 298920
rect 516600 298868 516652 298920
rect 517428 298868 517480 298920
rect 531228 298868 531280 298920
rect 538128 298868 538180 298920
rect 551560 298868 551612 298920
rect 557448 298868 557500 298920
rect 564532 298868 564584 298920
rect 565728 298868 565780 298920
rect 570144 298868 570196 298920
rect 472808 298800 472860 298852
rect 475384 298800 475436 298852
rect 480168 298800 480220 298852
rect 511724 298800 511776 298852
rect 513288 298800 513340 298852
rect 534448 298800 534500 298852
rect 535368 298800 535420 298852
rect 549904 298800 549956 298852
rect 551284 298800 551336 298852
rect 560484 298800 560536 298852
rect 7564 298732 7616 298784
rect 187240 298732 187292 298784
rect 214656 298732 214708 298784
rect 229376 298732 229428 298784
rect 230572 298732 230624 298784
rect 267556 298732 267608 298784
rect 268384 298732 268436 298784
rect 365720 298732 365772 298784
rect 367744 298732 367796 298784
rect 433892 298732 433944 298784
rect 438768 298732 438820 298784
rect 481732 298732 481784 298784
rect 482928 298732 482980 298784
rect 513380 298732 513432 298784
rect 516048 298732 516100 298784
rect 537760 298732 537812 298784
rect 539508 298732 539560 298784
rect 552296 298732 552348 298784
rect 567108 298732 567160 298784
rect 571800 298732 571852 298784
rect 582748 298775 582800 298784
rect 582748 298741 582757 298775
rect 582757 298741 582791 298775
rect 582791 298741 582800 298775
rect 582748 298732 582800 298741
rect 101404 298664 101456 298716
rect 248880 298664 248932 298716
rect 251732 298664 251784 298716
rect 262680 298664 262732 298716
rect 266360 298664 266412 298716
rect 278872 298664 278924 298716
rect 287796 298664 287848 298716
rect 315396 298664 315448 298716
rect 329104 298664 329156 298716
rect 394884 298664 394936 298716
rect 396724 298664 396776 298716
rect 453304 298664 453356 298716
rect 457352 298664 457404 298716
rect 460204 298664 460256 298716
rect 465540 298664 465592 298716
rect 466368 298664 466420 298716
rect 502064 298664 502116 298716
rect 509148 298664 509200 298716
rect 532056 298664 532108 298716
rect 114468 298596 114520 298648
rect 261024 298596 261076 298648
rect 274548 298596 274600 298648
rect 284576 298596 284628 298648
rect 298836 298596 298888 298648
rect 305828 298596 305880 298648
rect 310520 298596 310572 298648
rect 324964 298596 325016 298648
rect 121368 298528 121420 298580
rect 265900 298528 265952 298580
rect 278044 298528 278096 298580
rect 305644 298528 305696 298580
rect 360844 298528 360896 298580
rect 384304 298596 384356 298648
rect 387616 298596 387668 298648
rect 391204 298596 391256 298648
rect 392492 298596 392544 298648
rect 392584 298596 392636 298648
rect 397368 298596 397420 298648
rect 402244 298596 402296 298648
rect 458180 298596 458232 298648
rect 482284 298596 482336 298648
rect 507676 298596 507728 298648
rect 511908 298596 511960 298648
rect 533712 298664 533764 298716
rect 538864 298664 538916 298716
rect 548248 298664 548300 298716
rect 549168 298664 549220 298716
rect 558828 298664 558880 298716
rect 569316 298664 569368 298716
rect 570972 298664 571024 298716
rect 533344 298596 533396 298648
rect 540980 298596 541032 298648
rect 543096 298596 543148 298648
rect 553124 298596 553176 298648
rect 390008 298528 390060 298580
rect 87604 298460 87656 298512
rect 226984 298460 227036 298512
rect 250536 298460 250588 298512
rect 258816 298460 258868 298512
rect 338764 298460 338816 298512
rect 385224 298460 385276 298512
rect 386328 298460 386380 298512
rect 396816 298460 396868 298512
rect 83464 298392 83516 298444
rect 222108 298392 222160 298444
rect 317420 298392 317472 298444
rect 341340 298392 341392 298444
rect 345664 298392 345716 298444
rect 358728 298392 358780 298444
rect 387708 298392 387760 298444
rect 443276 298528 443328 298580
rect 444288 298528 444340 298580
rect 451188 298528 451240 298580
rect 492312 298528 492364 298580
rect 452568 298460 452620 298512
rect 458088 298460 458140 298512
rect 465724 298460 465776 298512
rect 489460 298460 489512 298512
rect 447692 298392 447744 298444
rect 474096 298392 474148 298444
rect 484216 298392 484268 298444
rect 487804 298392 487856 298444
rect 491944 298460 491996 298512
rect 499580 298528 499632 298580
rect 502984 298528 503036 298580
rect 497464 298460 497516 298512
rect 510160 298460 510212 298512
rect 521568 298528 521620 298580
rect 529204 298528 529256 298580
rect 542636 298528 542688 298580
rect 558828 298528 558880 298580
rect 566096 298528 566148 298580
rect 525524 298460 525576 298512
rect 536932 298460 536984 298512
rect 537484 298460 537536 298512
rect 545856 298460 545908 298512
rect 500868 298392 500920 298444
rect 508504 298392 508556 298444
rect 514208 298392 514260 298444
rect 520188 298392 520240 298444
rect 525064 298392 525116 298444
rect 532884 298392 532936 298444
rect 536104 298392 536156 298444
rect 544660 298392 544712 298444
rect 79324 298324 79376 298376
rect 217232 298324 217284 298376
rect 221464 298324 221516 298376
rect 288624 298324 288676 298376
rect 291016 298324 291068 298376
rect 338028 298324 338080 298376
rect 400128 298324 400180 298376
rect 411904 298324 411956 298376
rect 462228 298324 462280 298376
rect 483664 298324 483716 298376
rect 491208 298324 491260 298376
rect 496728 298324 496780 298376
rect 501604 298324 501656 298376
rect 510988 298324 511040 298376
rect 98644 298256 98696 298308
rect 231860 298256 231912 298308
rect 416044 298256 416096 298308
rect 424324 298256 424376 298308
rect 471980 298256 472032 298308
rect 480904 298256 480956 298308
rect 494704 298256 494756 298308
rect 500224 298256 500276 298308
rect 509332 298256 509384 298308
rect 511264 298256 511316 298308
rect 529572 298256 529624 298308
rect 561588 298256 561640 298308
rect 567752 298256 567804 298308
rect 105544 298188 105596 298240
rect 236736 298188 236788 298240
rect 406384 298188 406436 298240
rect 407120 298188 407172 298240
rect 423588 298188 423640 298240
rect 436008 298188 436060 298240
rect 447048 298188 447100 298240
rect 489000 298188 489052 298240
rect 233884 298120 233936 298172
rect 234528 298120 234580 298172
rect 263048 298120 263100 298172
rect 269120 298120 269172 298172
rect 448428 298120 448480 298172
rect 479524 298120 479576 298172
rect 480076 298120 480128 298172
rect 486424 298120 486476 298172
rect 498752 298188 498804 298240
rect 492036 298120 492088 298172
rect 504456 298188 504508 298240
rect 522304 298188 522356 298240
rect 528836 298188 528888 298240
rect 565084 298188 565136 298240
rect 569408 298188 569460 298240
rect 575388 298188 575440 298240
rect 577504 298188 577556 298240
rect 508228 298120 508280 298172
rect 518164 298120 518216 298172
rect 520648 298120 520700 298172
rect 554044 298120 554096 298172
rect 559656 298120 559708 298172
rect 566464 298120 566516 298172
rect 568580 298120 568632 298172
rect 576768 298120 576820 298172
rect 578332 298120 578384 298172
rect 140688 298052 140740 298104
rect 266360 298052 266412 298104
rect 341524 298052 341576 298104
rect 408684 298052 408736 298104
rect 413284 298052 413336 298104
rect 463884 298052 463936 298104
rect 135168 297984 135220 298036
rect 263692 297984 263744 298036
rect 267004 297984 267056 298036
rect 330024 297984 330076 298036
rect 343548 297984 343600 298036
rect 418436 297984 418488 298036
rect 418804 297984 418856 298036
rect 468760 297984 468812 298036
rect 133788 297916 133840 297968
rect 273996 297916 274048 297968
rect 323584 297916 323636 297968
rect 403808 297916 403860 297968
rect 407028 297916 407080 297968
rect 461492 297916 461544 297968
rect 489184 297916 489236 297968
rect 517060 297916 517112 297968
rect 129648 297848 129700 297900
rect 271604 297848 271656 297900
rect 305736 297848 305788 297900
rect 391664 297848 391716 297900
rect 111064 297780 111116 297832
rect 257804 297780 257856 297832
rect 260104 297780 260156 297832
rect 349436 297780 349488 297832
rect 360844 297780 360896 297832
rect 401416 297848 401468 297900
rect 403624 297848 403676 297900
rect 459008 297848 459060 297900
rect 461584 297848 461636 297900
rect 490656 297848 490708 297900
rect 400864 297780 400916 297832
rect 456616 297780 456668 297832
rect 468484 297780 468536 297832
rect 502800 297780 502852 297832
rect 104164 297712 104216 297764
rect 252928 297712 252980 297764
rect 280804 297712 280856 297764
rect 373816 297712 373868 297764
rect 395988 297712 396040 297764
rect 454132 297712 454184 297764
rect 471244 297712 471296 297764
rect 505284 297712 505336 297764
rect 93124 297644 93176 297696
rect 245660 297644 245712 297696
rect 268476 297644 268528 297696
rect 361672 297644 361724 297696
rect 392676 297644 392728 297696
rect 451740 297644 451792 297696
rect 464344 297644 464396 297696
rect 500408 297644 500460 297696
rect 88984 297576 89036 297628
rect 243176 297576 243228 297628
rect 269764 297576 269816 297628
rect 366548 297576 366600 297628
rect 389824 297576 389876 297628
rect 449256 297576 449308 297628
rect 457444 297576 457496 297628
rect 495532 297576 495584 297628
rect 86224 297508 86276 297560
rect 240784 297508 240836 297560
rect 271788 297508 271840 297560
rect 368940 297508 368992 297560
rect 382188 297508 382240 297560
rect 444380 297508 444432 297560
rect 453304 297508 453356 297560
rect 493140 297508 493192 297560
rect 495348 297508 495400 297560
rect 522028 297508 522080 297560
rect 57244 297440 57296 297492
rect 211528 297440 211580 297492
rect 244924 297440 244976 297492
rect 346676 297440 346728 297492
rect 378048 297440 378100 297492
rect 441988 297440 442040 297492
rect 447784 297440 447836 297492
rect 488264 297440 488316 297492
rect 491116 297440 491168 297492
rect 519912 297440 519964 297492
rect 14464 297372 14516 297424
rect 192116 297372 192168 297424
rect 242164 297372 242216 297424
rect 344652 297372 344704 297424
rect 350356 297372 350408 297424
rect 423312 297372 423364 297424
rect 425704 297372 425756 297424
rect 473636 297372 473688 297424
rect 484308 297372 484360 297424
rect 515036 297372 515088 297424
rect 179328 297304 179380 297356
rect 305276 297304 305328 297356
rect 320824 297304 320876 297356
rect 379520 297304 379572 297356
rect 414664 297304 414716 297356
rect 466276 297304 466328 297356
rect 144828 297236 144880 297288
rect 268844 297236 268896 297288
rect 356704 297236 356756 297288
rect 411168 297236 411220 297288
rect 428464 297236 428516 297288
rect 476028 297236 476080 297288
rect 142068 297168 142120 297220
rect 262864 297168 262916 297220
rect 264244 297168 264296 297220
rect 337292 297168 337344 297220
rect 370504 297168 370556 297220
rect 406292 297168 406344 297220
rect 432604 297168 432656 297220
rect 478512 297168 478564 297220
rect 246304 297100 246356 297152
rect 332416 297100 332468 297152
rect 447876 297100 447928 297152
rect 480628 297100 480680 297152
rect 250444 297032 250496 297084
rect 322664 297032 322716 297084
rect 453396 297032 453448 297084
rect 485780 297032 485832 297084
rect 258724 296964 258776 297016
rect 325148 296964 325200 297016
rect 262864 296896 262916 296948
rect 327540 296896 327592 296948
rect 177948 296624 178000 296676
rect 303712 296624 303764 296676
rect 309784 296624 309836 296676
rect 380992 296624 381044 296676
rect 158628 296556 158680 296608
rect 288624 296556 288676 296608
rect 318064 296556 318116 296608
rect 398932 296556 398984 296608
rect 147588 296488 147640 296540
rect 281356 296488 281408 296540
rect 287704 296488 287756 296540
rect 368480 296488 368532 296540
rect 151728 296420 151780 296472
rect 285772 296420 285824 296472
rect 304264 296420 304316 296472
rect 386512 296420 386564 296472
rect 113088 296352 113140 296404
rect 259552 296352 259604 296404
rect 273904 296352 273956 296404
rect 357532 296352 357584 296404
rect 108304 296284 108356 296336
rect 255412 296284 255464 296336
rect 298744 296284 298796 296336
rect 383660 296284 383712 296336
rect 99288 296216 99340 296268
rect 249800 296216 249852 296268
rect 286324 296216 286376 296268
rect 376852 296216 376904 296268
rect 95148 296148 95200 296200
rect 246948 296148 247000 296200
rect 262956 296148 263008 296200
rect 361580 296148 361632 296200
rect 376024 296148 376076 296200
rect 432052 296148 432104 296200
rect 54484 296080 54536 296132
rect 214012 296080 214064 296132
rect 240784 296080 240836 296132
rect 343640 296080 343692 296132
rect 370596 296080 370648 296132
rect 434812 296080 434864 296132
rect 47584 296012 47636 296064
rect 208400 296012 208452 296064
rect 223488 296012 223540 296064
rect 335452 296012 335504 296064
rect 375288 296012 375340 296064
rect 440332 296012 440384 296064
rect 25504 295944 25556 295996
rect 197452 295944 197504 295996
rect 209688 295944 209740 295996
rect 325792 295944 325844 295996
rect 336648 295944 336700 295996
rect 412732 295944 412784 295996
rect 439504 295944 439556 295996
rect 483112 295944 483164 295996
rect 148968 295876 149020 295928
rect 274548 295876 274600 295928
rect 291844 295876 291896 295928
rect 371332 295876 371384 295928
rect 256056 295808 256108 295860
rect 338212 295808 338264 295860
rect 251824 295740 251876 295792
rect 332600 295740 332652 295792
rect 124128 294856 124180 294908
rect 230572 294856 230624 294908
rect 117228 294788 117280 294840
rect 251732 294788 251784 294840
rect 119988 294720 120040 294772
rect 258080 294720 258132 294772
rect 51816 294652 51868 294704
rect 205732 294652 205784 294704
rect 32404 294584 32456 294636
rect 201592 294584 201644 294636
rect 231768 294584 231820 294636
rect 317420 294584 317472 294636
rect 3056 293904 3108 293956
rect 51724 293904 51776 293956
rect 582656 258927 582708 258936
rect 582656 258893 582665 258927
rect 582665 258893 582699 258927
rect 582699 258893 582708 258927
rect 582656 258884 582708 258893
rect 3148 255212 3200 255264
rect 40684 255212 40736 255264
rect 3516 241408 3568 241460
rect 39396 241408 39448 241460
rect 3056 202784 3108 202836
rect 137284 202784 137336 202836
rect 137928 202104 137980 202156
rect 276112 202104 276164 202156
rect 276664 202104 276716 202156
rect 367192 202104 367244 202156
rect 153108 188300 153160 188352
rect 285680 188300 285732 188352
rect 582564 165903 582616 165912
rect 582564 165869 582573 165903
rect 582573 165869 582607 165903
rect 582607 165869 582616 165903
rect 582564 165860 582616 165869
rect 3240 164160 3292 164212
rect 180064 164160 180116 164212
rect 582472 152711 582524 152720
rect 582472 152677 582481 152711
rect 582481 152677 582515 152711
rect 582515 152677 582524 152711
rect 582472 152668 582524 152677
rect 274088 141380 274140 141432
rect 340972 141380 341024 141432
rect 240968 140020 241020 140072
rect 320272 140020 320324 140072
rect 240876 139340 240928 139392
rect 579804 139340 579856 139392
rect 182916 113092 182968 113144
rect 579988 113092 580040 113144
rect 3424 111732 3476 111784
rect 15844 111732 15896 111784
rect 3424 97928 3476 97980
rect 36544 97928 36596 97980
rect 183008 86912 183060 86964
rect 580172 86912 580224 86964
rect 3148 85484 3200 85536
rect 39304 85484 39356 85536
rect 181904 73108 181956 73160
rect 580172 73108 580224 73160
rect 3424 71680 3476 71732
rect 22744 71680 22796 71732
rect 155868 48968 155920 49020
rect 288532 48968 288584 49020
rect 183100 46860 183152 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 61384 45500 61436 45552
rect 39304 39312 39356 39364
rect 204352 39312 204404 39364
rect 181996 33056 182048 33108
rect 579804 33056 579856 33108
rect 3424 20612 3476 20664
rect 583760 20612 583812 20664
rect 182088 20544 182140 20596
rect 580172 20544 580224 20596
rect 22744 19932 22796 19984
rect 194600 19932 194652 19984
rect 312636 18572 312688 18624
rect 396172 18572 396224 18624
rect 195888 17212 195940 17264
rect 316132 17212 316184 17264
rect 289084 14628 289136 14680
rect 374000 14628 374052 14680
rect 271144 14560 271196 14612
rect 358912 14560 358964 14612
rect 267096 14492 267148 14544
rect 364340 14492 364392 14544
rect 81348 14424 81400 14476
rect 237472 14424 237524 14476
rect 238024 14424 238076 14476
rect 339592 14424 339644 14476
rect 169668 13132 169720 13184
rect 250536 13132 250588 13184
rect 253388 13132 253440 13184
rect 334072 13132 334124 13184
rect 200028 13064 200080 13116
rect 312544 13064 312596 13116
rect 197268 12180 197320 12232
rect 273996 12180 274048 12232
rect 251088 12112 251140 12164
rect 353392 12112 353444 12164
rect 188988 12044 189040 12096
rect 300124 12044 300176 12096
rect 132408 11976 132460 12028
rect 253296 11976 253348 12028
rect 182088 11908 182140 11960
rect 306472 11908 306524 11960
rect 176568 11840 176620 11892
rect 302332 11840 302384 11892
rect 359464 11840 359516 11892
rect 427912 11840 427964 11892
rect 154212 11772 154264 11824
rect 288440 11772 288492 11824
rect 354588 11772 354640 11824
rect 425060 11772 425112 11824
rect 144736 11704 144788 11756
rect 281540 11704 281592 11756
rect 300768 11704 300820 11756
rect 389272 11704 389324 11756
rect 194508 10956 194560 11008
rect 287796 10956 287848 11008
rect 161296 10888 161348 10940
rect 258816 10888 258868 10940
rect 259368 10888 259420 10940
rect 358820 10888 358872 10940
rect 165528 10820 165580 10872
rect 253204 10820 253256 10872
rect 253848 10820 253900 10872
rect 356060 10820 356112 10872
rect 190368 10752 190420 10804
rect 296076 10752 296128 10804
rect 183468 10684 183520 10736
rect 298836 10684 298888 10736
rect 186136 10616 186188 10668
rect 305828 10616 305880 10668
rect 126888 10548 126940 10600
rect 263048 10548 263100 10600
rect 269856 10548 269908 10600
rect 352012 10548 352064 10600
rect 136456 10480 136508 10532
rect 276020 10480 276072 10532
rect 296628 10480 296680 10532
rect 385132 10480 385184 10532
rect 122748 10412 122800 10464
rect 266452 10412 266504 10464
rect 276756 10412 276808 10464
rect 371240 10412 371292 10464
rect 119804 10344 119856 10396
rect 263600 10344 263652 10396
rect 264888 10344 264940 10396
rect 363052 10344 363104 10396
rect 363604 10344 363656 10396
rect 430672 10344 430724 10396
rect 3424 10276 3476 10328
rect 172428 10208 172480 10260
rect 246396 10208 246448 10260
rect 156604 9596 156656 9648
rect 289912 9596 289964 9648
rect 149520 9528 149572 9580
rect 284392 9528 284444 9580
rect 153016 9460 153068 9512
rect 287060 9460 287112 9512
rect 145932 9392 145984 9444
rect 283012 9392 283064 9444
rect 142436 9324 142488 9376
rect 280252 9324 280304 9376
rect 138848 9256 138900 9308
rect 277400 9256 277452 9308
rect 135260 9188 135312 9240
rect 274732 9188 274784 9240
rect 115204 9120 115256 9172
rect 260932 9120 260984 9172
rect 108120 9052 108172 9104
rect 256700 9052 256752 9104
rect 111616 8984 111668 9036
rect 259460 8984 259512 9036
rect 104532 8916 104584 8968
rect 253940 8916 253992 8968
rect 160100 8848 160152 8900
rect 292672 8848 292724 8900
rect 206192 8780 206244 8832
rect 324320 8780 324372 8832
rect 213368 8712 213420 8764
rect 328460 8712 328512 8764
rect 209780 8644 209832 8696
rect 325700 8644 325752 8696
rect 216864 8576 216916 8628
rect 331220 8576 331272 8628
rect 220452 8508 220504 8560
rect 333980 8508 334032 8560
rect 227536 8440 227588 8492
rect 338120 8440 338172 8492
rect 223948 8372 224000 8424
rect 335360 8372 335412 8424
rect 73804 8236 73856 8288
rect 233332 8236 233384 8288
rect 70308 8168 70360 8220
rect 230480 8168 230532 8220
rect 66720 8100 66772 8152
rect 227812 8100 227864 8152
rect 63224 8032 63276 8084
rect 225052 8032 225104 8084
rect 59636 7964 59688 8016
rect 223672 7964 223724 8016
rect 56048 7896 56100 7948
rect 220912 7896 220964 7948
rect 251180 7896 251232 7948
rect 354772 7896 354824 7948
rect 52552 7828 52604 7880
rect 218152 7828 218204 7880
rect 247592 7828 247644 7880
rect 351920 7828 351972 7880
rect 48964 7760 49016 7812
rect 215392 7760 215444 7812
rect 244096 7760 244148 7812
rect 349160 7760 349212 7812
rect 44272 7692 44324 7744
rect 212540 7692 212592 7744
rect 240508 7692 240560 7744
rect 347872 7692 347924 7744
rect 40684 7624 40736 7676
rect 209872 7624 209924 7676
rect 233424 7624 233476 7676
rect 342260 7624 342312 7676
rect 37188 7556 37240 7608
rect 207112 7556 207164 7608
rect 237012 7556 237064 7608
rect 345112 7556 345164 7608
rect 371700 7556 371752 7608
rect 436744 7556 436796 7608
rect 77392 7488 77444 7540
rect 234712 7488 234764 7540
rect 101036 7420 101088 7472
rect 251272 7420 251324 7472
rect 128176 7352 128228 7404
rect 270500 7352 270552 7404
rect 158904 7284 158956 7336
rect 291200 7284 291252 7336
rect 163688 7216 163740 7268
rect 294052 7216 294104 7268
rect 167184 7148 167236 7200
rect 296812 7148 296864 7200
rect 170772 7080 170824 7132
rect 299572 7080 299624 7132
rect 174268 7012 174320 7064
rect 302240 7012 302292 7064
rect 162492 6808 162544 6860
rect 293960 6808 294012 6860
rect 130568 6740 130620 6792
rect 271972 6740 272024 6792
rect 374092 6740 374144 6792
rect 438860 6740 438912 6792
rect 126980 6672 127032 6724
rect 269212 6672 269264 6724
rect 370688 6672 370740 6724
rect 436192 6672 436244 6724
rect 97448 6604 97500 6656
rect 248512 6604 248564 6656
rect 367008 6604 367060 6656
rect 434720 6604 434772 6656
rect 93952 6536 94004 6588
rect 247132 6536 247184 6588
rect 339868 6536 339920 6588
rect 410524 6536 410576 6588
rect 90456 6468 90508 6520
rect 244280 6468 244332 6520
rect 292580 6468 292632 6520
rect 382372 6468 382424 6520
rect 86868 6400 86920 6452
rect 241612 6400 241664 6452
rect 288992 6400 289044 6452
rect 380900 6400 380952 6452
rect 389456 6400 389508 6452
rect 449164 6400 449216 6452
rect 83280 6332 83332 6384
rect 238852 6332 238904 6384
rect 285404 6332 285456 6384
rect 378140 6332 378192 6384
rect 382372 6332 382424 6384
rect 443644 6332 443696 6384
rect 79692 6264 79744 6316
rect 237380 6264 237432 6316
rect 281908 6264 281960 6316
rect 375472 6264 375524 6316
rect 384764 6264 384816 6316
rect 445852 6264 445904 6316
rect 8760 6196 8812 6248
rect 187792 6196 187844 6248
rect 190828 6196 190880 6248
rect 313372 6196 313424 6248
rect 346952 6196 347004 6248
rect 421012 6196 421064 6248
rect 4068 6128 4120 6180
rect 184940 6128 184992 6180
rect 187332 6128 187384 6180
rect 310612 6128 310664 6180
rect 311624 6128 311676 6180
rect 393412 6128 393464 6180
rect 501788 6128 501840 6180
rect 525156 6128 525208 6180
rect 166080 6060 166132 6112
rect 296720 6060 296772 6112
rect 169576 5992 169628 6044
rect 298192 5992 298244 6044
rect 173164 5924 173216 5976
rect 300860 5924 300912 5976
rect 176660 5856 176712 5908
rect 303620 5856 303672 5908
rect 180248 5788 180300 5840
rect 306380 5788 306432 5840
rect 183744 5720 183796 5772
rect 307852 5720 307904 5772
rect 194416 5652 194468 5704
rect 316040 5652 316092 5704
rect 197912 5584 197964 5636
rect 317512 5584 317564 5636
rect 47860 5448 47912 5500
rect 215300 5448 215352 5500
rect 306748 5448 306800 5500
rect 393320 5448 393372 5500
rect 33600 5380 33652 5432
rect 205640 5380 205692 5432
rect 303160 5380 303212 5432
rect 390560 5380 390612 5432
rect 30104 5312 30156 5364
rect 202880 5312 202932 5364
rect 299664 5312 299716 5364
rect 387800 5312 387852 5364
rect 26516 5244 26568 5296
rect 200212 5244 200264 5296
rect 231400 5244 231452 5296
rect 339500 5244 339552 5296
rect 342168 5244 342220 5296
rect 416872 5244 416924 5296
rect 17040 5176 17092 5228
rect 193312 5176 193364 5228
rect 215668 5176 215720 5228
rect 329840 5176 329892 5228
rect 335084 5176 335136 5228
rect 412640 5176 412692 5228
rect 21824 5108 21876 5160
rect 197360 5108 197412 5160
rect 212540 5108 212592 5160
rect 327080 5108 327132 5160
rect 331588 5108 331640 5160
rect 409880 5108 409932 5160
rect 12348 5040 12400 5092
rect 190552 5040 190604 5092
rect 201500 5040 201552 5092
rect 320180 5040 320232 5092
rect 320916 5040 320968 5092
rect 402980 5040 403032 5092
rect 7656 4972 7708 5024
rect 187700 4972 187752 5024
rect 205088 4972 205140 5024
rect 322940 4972 322992 5024
rect 324412 4972 324464 5024
rect 404452 4972 404504 5024
rect 2872 4904 2924 4956
rect 183560 4904 183612 4956
rect 202696 4904 202748 4956
rect 321560 4904 321612 4956
rect 328000 4904 328052 4956
rect 407212 4904 407264 4956
rect 572 4836 624 4888
rect 182180 4836 182232 4888
rect 192024 4836 192076 4888
rect 313280 4836 313332 4888
rect 313832 4836 313884 4888
rect 397460 4836 397512 4888
rect 459192 4836 459244 4888
rect 496912 4836 496964 4888
rect 1676 4768 1728 4820
rect 183652 4768 183704 4820
rect 184940 4768 184992 4820
rect 309140 4768 309192 4820
rect 310244 4768 310296 4820
rect 394792 4768 394844 4820
rect 420184 4768 420236 4820
rect 470600 4768 470652 4820
rect 51356 4700 51408 4752
rect 218060 4700 218112 4752
rect 317328 4700 317380 4752
rect 400220 4700 400272 4752
rect 54944 4632 54996 4684
rect 219532 4632 219584 4684
rect 338672 4632 338724 4684
rect 414112 4632 414164 4684
rect 62028 4564 62080 4616
rect 224960 4564 225012 4616
rect 345756 4564 345808 4616
rect 419540 4564 419592 4616
rect 58440 4496 58492 4548
rect 222200 4496 222252 4548
rect 349252 4496 349304 4548
rect 422300 4496 422352 4548
rect 65524 4428 65576 4480
rect 227720 4428 227772 4480
rect 352840 4428 352892 4480
rect 423772 4428 423824 4480
rect 72608 4360 72660 4412
rect 231952 4360 232004 4412
rect 356336 4360 356388 4412
rect 426532 4360 426584 4412
rect 69112 4292 69164 4344
rect 229192 4292 229244 4344
rect 359924 4292 359976 4344
rect 429200 4292 429252 4344
rect 76196 4224 76248 4276
rect 234620 4224 234672 4276
rect 363512 4224 363564 4276
rect 431960 4224 432012 4276
rect 67916 4088 67968 4140
rect 214656 4088 214708 4140
rect 226340 4088 226392 4140
rect 256056 4088 256108 4140
rect 258172 4088 258224 4140
rect 258724 4088 258776 4140
rect 259460 4088 259512 4140
rect 305460 4088 305512 4140
rect 319720 4088 319772 4140
rect 399484 4088 399536 4140
rect 402520 4088 402572 4140
rect 403532 4088 403584 4140
rect 463700 4088 463752 4140
rect 35164 4020 35216 4072
rect 38384 4020 38436 4072
rect 47584 4020 47636 4072
rect 57244 4020 57296 4072
rect 60832 4020 60884 4072
rect 221556 4020 221608 4072
rect 253388 4020 253440 4072
rect 257068 4020 257120 4072
rect 271144 4020 271196 4072
rect 298468 4020 298520 4072
rect 403624 4020 403676 4072
rect 459744 4020 459796 4072
rect 469220 4088 469272 4140
rect 469864 4088 469916 4140
rect 471244 4088 471296 4140
rect 468668 4020 468720 4072
rect 475752 4020 475804 4072
rect 505376 4088 505428 4140
rect 511172 4088 511224 4140
rect 500224 4020 500276 4072
rect 524236 4020 524288 4072
rect 529204 4020 529256 4072
rect 14740 3952 14792 4004
rect 18604 3952 18656 4004
rect 34796 3952 34848 4004
rect 51816 3952 51868 4004
rect 53748 3952 53800 4004
rect 210424 3952 210476 4004
rect 219256 3952 219308 4004
rect 251824 3952 251876 4004
rect 254676 3952 254728 4004
rect 273904 3952 273956 4004
rect 276020 3952 276072 4004
rect 291844 3952 291896 4004
rect 293684 3952 293736 4004
rect 298744 3952 298796 4004
rect 305552 3952 305604 4004
rect 391204 3952 391256 4004
rect 393044 3952 393096 4004
rect 396816 3952 396868 4004
rect 397736 3952 397788 4004
rect 455420 3952 455472 4004
rect 460388 3952 460440 4004
rect 486332 3952 486384 4004
rect 25320 3884 25372 3936
rect 29644 3884 29696 3936
rect 31300 3884 31352 3936
rect 39304 3884 39356 3936
rect 43076 3884 43128 3936
rect 211804 3884 211856 3936
rect 225144 3884 225196 3936
rect 264244 3884 264296 3936
rect 266544 3884 266596 3936
rect 268384 3884 268436 3936
rect 272432 3884 272484 3936
rect 279516 3884 279568 3936
rect 289084 3884 289136 3936
rect 382280 3884 382332 3936
rect 392584 3884 392636 3936
rect 454040 3884 454092 3936
rect 454500 3884 454552 3936
rect 480904 3884 480956 3936
rect 492036 3884 492088 3936
rect 504180 3884 504232 3936
rect 522304 3884 522356 3936
rect 24216 3816 24268 3868
rect 28908 3816 28960 3868
rect 27712 3748 27764 3800
rect 32404 3748 32456 3800
rect 35992 3816 36044 3868
rect 207020 3816 207072 3868
rect 234620 3816 234672 3868
rect 240784 3816 240836 3868
rect 274088 3816 274140 3868
rect 284300 3816 284352 3868
rect 376760 3816 376812 3868
rect 384304 3816 384356 3868
rect 390652 3816 390704 3868
rect 449992 3816 450044 3868
rect 461584 3816 461636 3868
rect 491944 3816 491996 3868
rect 497096 3816 497148 3868
rect 519452 3816 519504 3868
rect 531320 3816 531372 3868
rect 546684 3816 546736 3868
rect 20628 3680 20680 3732
rect 195980 3680 196032 3732
rect 211160 3748 211212 3800
rect 214472 3748 214524 3800
rect 201592 3680 201644 3732
rect 210976 3680 211028 3732
rect 262864 3748 262916 3800
rect 270040 3748 270092 3800
rect 263048 3680 263100 3732
rect 19432 3612 19484 3664
rect 196072 3612 196124 3664
rect 207388 3612 207440 3664
rect 258172 3612 258224 3664
rect 258264 3612 258316 3664
rect 259368 3612 259420 3664
rect 261760 3612 261812 3664
rect 262956 3612 263008 3664
rect 264152 3612 264204 3664
rect 264888 3612 264940 3664
rect 265348 3612 265400 3664
rect 267096 3612 267148 3664
rect 267740 3680 267792 3732
rect 269764 3680 269816 3732
rect 271236 3680 271288 3732
rect 271788 3680 271840 3732
rect 277124 3748 277176 3800
rect 371884 3748 371936 3800
rect 378876 3748 378928 3800
rect 380164 3748 380216 3800
rect 383568 3748 383620 3800
rect 432052 3748 432104 3800
rect 367100 3680 367152 3732
rect 369400 3680 369452 3732
rect 355232 3612 355284 3664
rect 365812 3612 365864 3664
rect 367744 3612 367796 3664
rect 368204 3612 368256 3664
rect 370596 3612 370648 3664
rect 372896 3680 372948 3732
rect 373908 3680 373960 3732
rect 379980 3680 380032 3732
rect 380808 3680 380860 3732
rect 381176 3680 381228 3732
rect 382188 3680 382240 3732
rect 11152 3544 11204 3596
rect 203892 3544 203944 3596
rect 13544 3476 13596 3528
rect 14464 3476 14516 3528
rect 5264 3408 5316 3460
rect 6460 3272 6512 3324
rect 7564 3272 7616 3324
rect 9956 3340 10008 3392
rect 181444 3476 181496 3528
rect 182088 3476 182140 3528
rect 182548 3476 182600 3528
rect 183468 3476 183520 3528
rect 188528 3476 188580 3528
rect 188988 3476 189040 3528
rect 190460 3476 190512 3528
rect 193220 3476 193272 3528
rect 194508 3476 194560 3528
rect 196808 3476 196860 3528
rect 197268 3476 197320 3528
rect 208584 3476 208636 3528
rect 209688 3476 209740 3528
rect 218060 3476 218112 3528
rect 246304 3476 246356 3528
rect 248788 3544 248840 3596
rect 249892 3476 249944 3528
rect 249984 3476 250036 3528
rect 251088 3476 251140 3528
rect 255872 3544 255924 3596
rect 357440 3544 357492 3596
rect 353484 3476 353536 3528
rect 354036 3476 354088 3528
rect 354588 3476 354640 3528
rect 362224 3544 362276 3596
rect 362316 3544 362368 3596
rect 430580 3544 430632 3596
rect 430856 3544 430908 3596
rect 432604 3544 432656 3596
rect 361120 3476 361172 3528
rect 363604 3476 363656 3528
rect 422576 3476 422628 3528
rect 423588 3476 423640 3528
rect 423772 3476 423824 3528
rect 425704 3476 425756 3528
rect 427268 3476 427320 3528
rect 428464 3476 428516 3528
rect 429660 3476 429712 3528
rect 430488 3476 430540 3528
rect 440240 3680 440292 3732
rect 433248 3612 433300 3664
rect 437940 3544 437992 3596
rect 439504 3544 439556 3596
rect 435364 3476 435416 3528
rect 435548 3476 435600 3528
rect 436008 3476 436060 3528
rect 436744 3476 436796 3528
rect 438124 3476 438176 3528
rect 441528 3748 441580 3800
rect 445024 3748 445076 3800
rect 447784 3748 447836 3800
rect 446220 3680 446272 3732
rect 447048 3680 447100 3732
rect 447416 3680 447468 3732
rect 465724 3748 465776 3800
rect 472256 3748 472308 3800
rect 504364 3748 504416 3800
rect 518164 3748 518216 3800
rect 521844 3748 521896 3800
rect 533344 3748 533396 3800
rect 456064 3680 456116 3732
rect 456892 3680 456944 3732
rect 493324 3680 493376 3732
rect 499396 3680 499448 3732
rect 502984 3680 503036 3732
rect 507676 3680 507728 3732
rect 529296 3680 529348 3732
rect 440424 3612 440476 3664
rect 479524 3612 479576 3664
rect 492312 3612 492364 3664
rect 474004 3544 474056 3596
rect 487804 3544 487856 3596
rect 488816 3544 488868 3596
rect 489828 3544 489880 3596
rect 489920 3544 489972 3596
rect 491208 3544 491260 3596
rect 493508 3544 493560 3596
rect 493968 3544 494020 3596
rect 495900 3544 495952 3596
rect 496728 3544 496780 3596
rect 498200 3612 498252 3664
rect 522396 3612 522448 3664
rect 536196 3680 536248 3732
rect 546684 3680 546736 3732
rect 548524 3680 548576 3732
rect 510068 3544 510120 3596
rect 525064 3544 525116 3596
rect 525432 3544 525484 3596
rect 543188 3612 543240 3664
rect 544384 3612 544436 3664
rect 471060 3476 471112 3528
rect 478052 3476 478104 3528
rect 479340 3476 479392 3528
rect 480168 3476 480220 3528
rect 482836 3476 482888 3528
rect 186412 3408 186464 3460
rect 189724 3408 189776 3460
rect 190368 3408 190420 3460
rect 199108 3408 199160 3460
rect 200028 3408 200080 3460
rect 200304 3408 200356 3460
rect 231032 3408 231084 3460
rect 231768 3408 231820 3460
rect 232228 3408 232280 3460
rect 241704 3408 241756 3460
rect 344560 3408 344612 3460
rect 345664 3408 345716 3460
rect 348056 3408 348108 3460
rect 413100 3408 413152 3460
rect 414664 3408 414716 3460
rect 415492 3408 415544 3460
rect 416688 3408 416740 3460
rect 421380 3408 421432 3460
rect 424324 3408 424376 3460
rect 426164 3408 426216 3460
rect 474740 3408 474792 3460
rect 15936 3340 15988 3392
rect 17224 3340 17276 3392
rect 32404 3340 32456 3392
rect 33784 3340 33836 3392
rect 39580 3340 39632 3392
rect 43444 3340 43496 3392
rect 45468 3340 45520 3392
rect 54484 3340 54536 3392
rect 75000 3340 75052 3392
rect 214564 3340 214616 3392
rect 222752 3340 222804 3392
rect 223488 3340 223540 3392
rect 238116 3340 238168 3392
rect 249064 3340 249116 3392
rect 252376 3340 252428 3392
rect 278044 3340 278096 3392
rect 278320 3340 278372 3392
rect 280804 3340 280856 3392
rect 283104 3340 283156 3392
rect 286324 3340 286376 3392
rect 286600 3340 286652 3392
rect 320824 3340 320876 3392
rect 322112 3340 322164 3392
rect 323584 3340 323636 3392
rect 330392 3340 330444 3392
rect 331864 3340 331916 3392
rect 41880 3272 41932 3324
rect 50160 3272 50212 3324
rect 79324 3272 79376 3324
rect 80888 3272 80940 3324
rect 81348 3272 81400 3324
rect 84476 3272 84528 3324
rect 86224 3272 86276 3324
rect 87972 3272 88024 3324
rect 88984 3272 89036 3324
rect 89168 3272 89220 3324
rect 90364 3272 90416 3324
rect 91560 3272 91612 3324
rect 93124 3272 93176 3324
rect 217324 3272 217376 3324
rect 228732 3272 228784 3324
rect 238024 3272 238076 3324
rect 18236 3204 18288 3256
rect 22744 3204 22796 3256
rect 23020 3204 23072 3256
rect 25504 3204 25556 3256
rect 57244 3204 57296 3256
rect 83464 3204 83516 3256
rect 85672 3204 85724 3256
rect 220084 3204 220136 3256
rect 235816 3204 235868 3256
rect 242164 3272 242216 3324
rect 246396 3272 246448 3324
rect 269856 3272 269908 3324
rect 274824 3272 274876 3324
rect 276756 3272 276808 3324
rect 287704 3272 287756 3324
rect 290188 3272 290240 3324
rect 309784 3272 309836 3324
rect 311440 3272 311492 3324
rect 312636 3272 312688 3324
rect 312728 3272 312780 3324
rect 326804 3272 326856 3324
rect 64328 3136 64380 3188
rect 87604 3136 87656 3188
rect 92756 3136 92808 3188
rect 221464 3136 221516 3188
rect 240968 3204 241020 3256
rect 242900 3204 242952 3256
rect 260104 3204 260156 3256
rect 260656 3204 260708 3256
rect 268476 3204 268528 3256
rect 273628 3204 273680 3256
rect 282184 3204 282236 3256
rect 291384 3204 291436 3256
rect 297272 3204 297324 3256
rect 304264 3204 304316 3256
rect 304356 3204 304408 3256
rect 305736 3204 305788 3256
rect 239312 3136 239364 3188
rect 244924 3136 244976 3188
rect 245200 3136 245252 3188
rect 255964 3136 256016 3188
rect 267004 3136 267056 3188
rect 294880 3136 294932 3188
rect 71504 3068 71556 3120
rect 98552 3068 98604 3120
rect 98644 3068 98696 3120
rect 99288 3068 99340 3120
rect 102232 3068 102284 3120
rect 104164 3068 104216 3120
rect 106924 3068 106976 3120
rect 107568 3068 107620 3120
rect 109316 3068 109368 3120
rect 111064 3068 111116 3120
rect 46664 3000 46716 3052
rect 50344 3000 50396 3052
rect 78588 3000 78640 3052
rect 82084 2932 82136 2984
rect 99840 3000 99892 3052
rect 224224 3068 224276 3120
rect 268844 3068 268896 3120
rect 276664 3068 276716 3120
rect 280712 3068 280764 3120
rect 284944 3068 284996 3120
rect 287796 3068 287848 3120
rect 295984 3068 296036 3120
rect 96252 2932 96304 2984
rect 101404 2932 101456 2984
rect 105728 2932 105780 2984
rect 108304 2932 108356 2984
rect 110512 2932 110564 2984
rect 226984 3000 227036 3052
rect 296076 3000 296128 3052
rect 296628 3000 296680 3052
rect 301964 3068 302016 3120
rect 316224 3204 316276 3256
rect 322204 3204 322256 3256
rect 323308 3204 323360 3256
rect 327724 3204 327776 3256
rect 391848 3272 391900 3324
rect 392676 3272 392728 3324
rect 395344 3272 395396 3324
rect 395988 3272 396040 3324
rect 398932 3272 398984 3324
rect 400864 3272 400916 3324
rect 401324 3272 401376 3324
rect 402244 3272 402296 3324
rect 406016 3340 406068 3392
rect 407028 3340 407080 3392
rect 407212 3340 407264 3392
rect 411904 3340 411956 3392
rect 414296 3340 414348 3392
rect 416044 3340 416096 3392
rect 404820 3272 404872 3324
rect 452108 3272 452160 3324
rect 453304 3272 453356 3324
rect 455696 3272 455748 3324
rect 457444 3272 457496 3324
rect 406384 3204 406436 3256
rect 410800 3204 410852 3256
rect 416688 3204 416740 3256
rect 418804 3204 418856 3256
rect 418988 3204 419040 3256
rect 462780 3340 462832 3392
rect 464344 3340 464396 3392
rect 465172 3340 465224 3392
rect 466368 3340 466420 3392
rect 478236 3408 478288 3460
rect 481732 3408 481784 3460
rect 482928 3408 482980 3460
rect 485228 3476 485280 3528
rect 485688 3476 485740 3528
rect 487620 3476 487672 3528
rect 489184 3476 489236 3528
rect 502984 3476 503036 3528
rect 503628 3476 503680 3528
rect 506480 3476 506532 3528
rect 507768 3476 507820 3528
rect 511264 3476 511316 3528
rect 511908 3476 511960 3528
rect 512460 3476 512512 3528
rect 513288 3476 513340 3528
rect 513564 3476 513616 3528
rect 515404 3476 515456 3528
rect 518348 3476 518400 3528
rect 518808 3476 518860 3528
rect 519544 3476 519596 3528
rect 520188 3476 520240 3528
rect 520740 3476 520792 3528
rect 521568 3476 521620 3528
rect 523040 3476 523092 3528
rect 526444 3476 526496 3528
rect 526628 3476 526680 3528
rect 527088 3476 527140 3528
rect 527824 3476 527876 3528
rect 536104 3544 536156 3596
rect 549076 3544 549128 3596
rect 554044 3544 554096 3596
rect 565636 3544 565688 3596
rect 569316 3544 569368 3596
rect 534908 3476 534960 3528
rect 535368 3476 535420 3528
rect 537208 3476 537260 3528
rect 538128 3476 538180 3528
rect 538404 3476 538456 3528
rect 539508 3476 539560 3528
rect 541992 3476 542044 3528
rect 543004 3476 543056 3528
rect 544384 3476 544436 3528
rect 545028 3476 545080 3528
rect 545488 3476 545540 3528
rect 547144 3476 547196 3528
rect 547880 3476 547932 3528
rect 549168 3476 549220 3528
rect 550272 3476 550324 3528
rect 551284 3476 551336 3528
rect 551468 3476 551520 3528
rect 551928 3476 551980 3528
rect 556160 3476 556212 3528
rect 557448 3476 557500 3528
rect 560852 3476 560904 3528
rect 561588 3476 561640 3528
rect 564440 3476 564492 3528
rect 565728 3476 565780 3528
rect 568028 3476 568080 3528
rect 569224 3476 569276 3528
rect 571524 3476 571576 3528
rect 572628 3476 572680 3528
rect 573916 3476 573968 3528
rect 575572 3476 575624 3528
rect 576308 3476 576360 3528
rect 576768 3476 576820 3528
rect 577412 3476 577464 3528
rect 578424 3476 578476 3528
rect 512092 3408 512144 3460
rect 514760 3408 514812 3460
rect 530584 3408 530636 3460
rect 554964 3408 555016 3460
rect 556804 3408 556856 3460
rect 559748 3408 559800 3460
rect 560944 3408 560996 3460
rect 570328 3408 570380 3460
rect 574192 3408 574244 3460
rect 478144 3340 478196 3392
rect 501604 3340 501656 3392
rect 508504 3340 508556 3392
rect 530124 3340 530176 3392
rect 531228 3340 531280 3392
rect 536104 3340 536156 3392
rect 540244 3340 540296 3392
rect 553768 3340 553820 3392
rect 561864 3340 561916 3392
rect 466276 3272 466328 3324
rect 468484 3272 468536 3324
rect 476948 3272 477000 3324
rect 497464 3272 497516 3324
rect 529020 3272 529072 3324
rect 537484 3272 537536 3324
rect 562048 3272 562100 3324
rect 566464 3272 566516 3324
rect 469312 3204 469364 3256
rect 474556 3204 474608 3256
rect 480536 3204 480588 3256
rect 569132 3204 569184 3256
rect 572904 3204 572956 3256
rect 338764 3136 338816 3188
rect 340972 3136 341024 3188
rect 416780 3136 416832 3188
rect 426440 3136 426492 3188
rect 428464 3136 428516 3188
rect 472624 3136 472676 3188
rect 473452 3136 473504 3188
rect 482284 3136 482336 3188
rect 532516 3136 532568 3188
rect 538864 3136 538916 3188
rect 539600 3136 539652 3188
rect 543096 3136 543148 3188
rect 552664 3136 552716 3188
rect 555424 3136 555476 3188
rect 563244 3136 563296 3188
rect 565084 3136 565136 3188
rect 583392 3136 583444 3188
rect 307944 3068 307996 3120
rect 311624 3068 311676 3120
rect 324964 3068 325016 3120
rect 325608 3068 325660 3120
rect 370504 3068 370556 3120
rect 376484 3068 376536 3120
rect 394240 3068 394292 3120
rect 396724 3068 396776 3120
rect 411260 3068 411312 3120
rect 411904 3068 411956 3120
rect 460204 3068 460256 3120
rect 463976 3068 464028 3120
rect 483664 3068 483716 3120
rect 318524 3000 318576 3052
rect 360844 3000 360896 3052
rect 387156 3000 387208 3052
rect 387708 3000 387760 3052
rect 396540 3000 396592 3052
rect 409604 3000 409656 3052
rect 413284 3000 413336 3052
rect 417884 3000 417936 3052
rect 439136 3000 439188 3052
rect 474096 3000 474148 3052
rect 486424 3000 486476 3052
rect 487068 3000 487120 3052
rect 494704 3000 494756 3052
rect 495348 3000 495400 3052
rect 578608 3000 578660 3052
rect 579620 3000 579672 3052
rect 114008 2932 114060 2984
rect 114468 2932 114520 2984
rect 116400 2932 116452 2984
rect 117228 2932 117280 2984
rect 118792 2932 118844 2984
rect 119804 2932 119856 2984
rect 122288 2932 122340 2984
rect 122748 2932 122800 2984
rect 123484 2932 123536 2984
rect 124128 2932 124180 2984
rect 125876 2932 125928 2984
rect 126888 2932 126940 2984
rect 105544 2864 105596 2916
rect 117596 2864 117648 2916
rect 232504 2932 232556 2984
rect 309048 2932 309100 2984
rect 329104 2932 329156 2984
rect 332692 2932 332744 2984
rect 356704 2932 356756 2984
rect 357532 2932 357584 2984
rect 359464 2932 359516 2984
rect 364616 2932 364668 2984
rect 376024 2932 376076 2984
rect 420920 2932 420972 2984
rect 442264 2932 442316 2984
rect 442632 2932 442684 2984
rect 476764 2932 476816 2984
rect 557356 2932 557408 2984
rect 558184 2932 558236 2984
rect 124680 2796 124732 2848
rect 233884 2864 233936 2916
rect 315028 2864 315080 2916
rect 318064 2864 318116 2916
rect 329196 2864 329248 2916
rect 131764 2796 131816 2848
rect 132408 2796 132460 2848
rect 132960 2796 133012 2848
rect 133788 2796 133840 2848
rect 134156 2796 134208 2848
rect 135168 2796 135220 2848
rect 140044 2796 140096 2848
rect 140688 2796 140740 2848
rect 141240 2796 141292 2848
rect 142068 2796 142120 2848
rect 143540 2796 143592 2848
rect 144828 2796 144880 2848
rect 147128 2796 147180 2848
rect 147588 2796 147640 2848
rect 148324 2796 148376 2848
rect 148968 2796 149020 2848
rect 150624 2796 150676 2848
rect 151728 2796 151780 2848
rect 151820 2796 151872 2848
rect 153108 2796 153160 2848
rect 155408 2796 155460 2848
rect 155868 2796 155920 2848
rect 157800 2796 157852 2848
rect 158628 2796 158680 2848
rect 164884 2796 164936 2848
rect 165528 2796 165580 2848
rect 168380 2796 168432 2848
rect 169668 2796 169720 2848
rect 171968 2796 172020 2848
rect 172428 2796 172480 2848
rect 175464 2796 175516 2848
rect 176568 2796 176620 2848
rect 189172 2796 189224 2848
rect 229836 2796 229888 2848
rect 231400 2796 231452 2848
rect 333888 2796 333940 2848
rect 347044 2864 347096 2916
rect 388260 2864 388312 2916
rect 389824 2864 389876 2916
rect 453212 2864 453264 2916
rect 453304 2864 453356 2916
rect 475384 2864 475436 2916
rect 572720 2864 572772 2916
rect 574008 2864 574060 2916
rect 341524 2796 341576 2848
rect 434444 2796 434496 2848
rect 447876 2796 447928 2848
rect 448612 2796 448664 2848
rect 461492 2796 461544 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 15844 703792 15896 703798
rect 15844 703734 15896 703740
rect 3422 700360 3478 700369
rect 3422 700295 3478 700304
rect 3056 672036 3108 672042
rect 3056 671978 3108 671984
rect 3068 671265 3096 671978
rect 3054 671256 3110 671265
rect 3054 671191 3110 671200
rect 3240 633412 3292 633418
rect 3240 633354 3292 633360
rect 3252 632097 3280 633354
rect 3238 632088 3294 632097
rect 3238 632023 3294 632032
rect 3332 619608 3384 619614
rect 3332 619550 3384 619556
rect 3344 619177 3372 619550
rect 3330 619168 3386 619177
rect 3330 619103 3386 619112
rect 3240 607164 3292 607170
rect 3240 607106 3292 607112
rect 3252 606121 3280 607106
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3148 580984 3200 580990
rect 3148 580926 3200 580932
rect 3160 580009 3188 580926
rect 3146 580000 3202 580009
rect 3146 579935 3202 579944
rect 2872 528556 2924 528562
rect 2872 528498 2924 528504
rect 2884 527921 2912 528498
rect 2870 527912 2926 527921
rect 2870 527847 2926 527856
rect 3240 463684 3292 463690
rect 3240 463626 3292 463632
rect 3252 462641 3280 463626
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3240 398812 3292 398818
rect 3240 398754 3292 398760
rect 3252 397497 3280 398754
rect 3238 397488 3294 397497
rect 3238 397423 3294 397432
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 3068 293185 3096 293898
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3436 188873 3464 700295
rect 8128 699990 8156 703520
rect 14464 702296 14516 702302
rect 14464 702238 14516 702244
rect 8116 699984 8168 699990
rect 8116 699926 8168 699932
rect 3516 684480 3568 684486
rect 3516 684422 3568 684428
rect 3528 684321 3556 684422
rect 3514 684312 3570 684321
rect 3514 684247 3570 684256
rect 3516 658232 3568 658238
rect 3514 658200 3516 658209
rect 3568 658200 3570 658209
rect 3514 658135 3570 658144
rect 3516 567180 3568 567186
rect 3516 567122 3568 567128
rect 3528 566953 3556 567122
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3516 554736 3568 554742
rect 3516 554678 3568 554684
rect 3528 553897 3556 554678
rect 3514 553888 3570 553897
rect 3514 553823 3570 553832
rect 3516 516112 3568 516118
rect 3516 516054 3568 516060
rect 3528 514865 3556 516054
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 14476 502314 14504 702238
rect 14556 699780 14608 699786
rect 14556 699722 14608 699728
rect 14568 658238 14596 699722
rect 14556 658232 14608 658238
rect 14556 658174 14608 658180
rect 3516 502308 3568 502314
rect 3516 502250 3568 502256
rect 14464 502308 14516 502314
rect 14464 502250 14516 502256
rect 3528 501809 3556 502250
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 3516 476060 3568 476066
rect 3516 476002 3568 476008
rect 3528 475697 3556 476002
rect 3514 475688 3570 475697
rect 3514 475623 3570 475632
rect 3516 423632 3568 423638
rect 3514 423600 3516 423609
rect 3568 423600 3570 423609
rect 3514 423535 3570 423544
rect 3516 372564 3568 372570
rect 3516 372506 3568 372512
rect 3528 371385 3556 372506
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 7564 298784 7616 298790
rect 7564 298726 7616 298732
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3422 138000 3478 138009
rect 3422 137935 3478 137944
rect 3436 136785 3464 137935
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3330 59256 3386 59265
rect 3330 59191 3386 59200
rect 3344 58585 3372 59191
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3330 33144 3386 33153
rect 3330 33079 3386 33088
rect 3344 32473 3372 33079
rect 3330 32464 3386 32473
rect 3330 32399 3386 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 10328 3476 10334
rect 3424 10270 3476 10276
rect 3436 6497 3464 10270
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 4898
rect 4080 480 4108 6122
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 7576 3330 7604 298726
rect 14464 297424 14516 297430
rect 14464 297366 14516 297372
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 6460 3324 6512 3330
rect 6460 3266 6512 3272
rect 7564 3324 7616 3330
rect 7564 3266 7616 3272
rect 6472 480 6500 3266
rect 7668 480 7696 4966
rect 8772 480 8800 6190
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9968 480 9996 3334
rect 11164 480 11192 3538
rect 12360 480 12388 5034
rect 14476 3534 14504 297366
rect 15856 111790 15884 703734
rect 22744 703724 22796 703730
rect 22744 703666 22796 703672
rect 18604 702364 18656 702370
rect 18604 702306 18656 702312
rect 17222 701584 17278 701593
rect 17222 701519 17278 701528
rect 17236 398818 17264 701519
rect 18616 516118 18644 702306
rect 18696 699848 18748 699854
rect 18696 699790 18748 699796
rect 18708 672042 18736 699790
rect 18696 672036 18748 672042
rect 18696 671978 18748 671984
rect 18604 516112 18656 516118
rect 18604 516054 18656 516060
rect 17224 398812 17276 398818
rect 17224 398754 17276 398760
rect 18604 298920 18656 298926
rect 18604 298862 18656 298868
rect 17224 298852 17276 298858
rect 17224 298794 17276 298800
rect 15844 111784 15896 111790
rect 15844 111726 15896 111732
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 13556 480 13584 3470
rect 14752 480 14780 3946
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15948 480 15976 3334
rect 17052 480 17080 5170
rect 17236 3398 17264 298794
rect 18616 4010 18644 298862
rect 22756 71738 22784 703666
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 235446 703760 235502 703769
rect 235446 703695 235502 703704
rect 235460 703610 235488 703695
rect 235368 703582 235488 703610
rect 24320 700194 24348 703520
rect 35164 702432 35216 702438
rect 35164 702374 35216 702380
rect 25502 701720 25558 701729
rect 25502 701655 25558 701664
rect 24308 700188 24360 700194
rect 24308 700130 24360 700136
rect 25516 411262 25544 701655
rect 29642 701448 29698 701457
rect 29642 701383 29698 701392
rect 25504 411256 25556 411262
rect 25504 411198 25556 411204
rect 29656 358766 29684 701383
rect 33782 701312 33838 701321
rect 32404 701276 32456 701282
rect 33782 701247 33838 701256
rect 32404 701218 32456 701224
rect 32416 449886 32444 701218
rect 32496 700120 32548 700126
rect 32496 700062 32548 700068
rect 32508 607170 32536 700062
rect 32496 607164 32548 607170
rect 32496 607106 32548 607112
rect 32404 449880 32456 449886
rect 32404 449822 32456 449828
rect 29644 358760 29696 358766
rect 29644 358702 29696 358708
rect 33796 306338 33824 701247
rect 33876 699712 33928 699718
rect 33876 699654 33928 699660
rect 33888 554742 33916 699654
rect 33876 554736 33928 554742
rect 33876 554678 33928 554684
rect 35176 463690 35204 702374
rect 39304 701344 39356 701350
rect 39304 701286 39356 701292
rect 36544 700528 36596 700534
rect 36544 700470 36596 700476
rect 35256 700052 35308 700058
rect 35256 699994 35308 700000
rect 35268 619614 35296 699994
rect 35256 619608 35308 619614
rect 35256 619550 35308 619556
rect 35164 463684 35216 463690
rect 35164 463626 35216 463632
rect 33784 306332 33836 306338
rect 33784 306274 33836 306280
rect 35164 299192 35216 299198
rect 35164 299134 35216 299140
rect 33784 299056 33836 299062
rect 33784 298998 33836 299004
rect 29644 298988 29696 298994
rect 29644 298930 29696 298936
rect 25504 295996 25556 296002
rect 25504 295938 25556 295944
rect 22744 71732 22796 71738
rect 22744 71674 22796 71680
rect 22744 19984 22796 19990
rect 22744 19926 22796 19932
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 18236 3256 18288 3262
rect 18236 3198 18288 3204
rect 18248 480 18276 3198
rect 19444 480 19472 3606
rect 20640 480 20668 3674
rect 21836 480 21864 5102
rect 22756 3262 22784 19926
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 24216 3868 24268 3874
rect 24216 3810 24268 3816
rect 22744 3256 22796 3262
rect 22744 3198 22796 3204
rect 23020 3256 23072 3262
rect 23020 3198 23072 3204
rect 23032 480 23060 3198
rect 24228 480 24256 3810
rect 25332 480 25360 3878
rect 25516 3262 25544 295938
rect 26516 5296 26568 5302
rect 26516 5238 26568 5244
rect 25504 3256 25556 3262
rect 25504 3198 25556 3204
rect 26528 480 26556 5238
rect 29656 3942 29684 298930
rect 32404 294636 32456 294642
rect 32404 294578 32456 294584
rect 30104 5364 30156 5370
rect 30104 5306 30156 5312
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 28908 3868 28960 3874
rect 28908 3810 28960 3816
rect 27712 3800 27764 3806
rect 27712 3742 27764 3748
rect 27724 480 27752 3742
rect 28920 480 28948 3810
rect 30116 480 30144 5306
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 31312 480 31340 3878
rect 32416 3806 32444 294578
rect 33600 5432 33652 5438
rect 33600 5374 33652 5380
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 32416 480 32444 3334
rect 33612 480 33640 5374
rect 33796 3398 33824 298998
rect 35176 4078 35204 299134
rect 36556 97986 36584 700470
rect 36544 97980 36596 97986
rect 36544 97922 36596 97928
rect 39316 85542 39344 701286
rect 39394 701176 39450 701185
rect 39394 701111 39450 701120
rect 39408 241466 39436 701111
rect 40512 701049 40540 703520
rect 51722 701856 51778 701865
rect 51722 701791 51778 701800
rect 40498 701040 40554 701049
rect 40498 700975 40554 700984
rect 40776 699916 40828 699922
rect 40776 699858 40828 699864
rect 40682 699816 40738 699825
rect 40682 699751 40738 699760
rect 40696 255270 40724 699751
rect 40788 567186 40816 699858
rect 40776 567180 40828 567186
rect 40776 567122 40828 567128
rect 50344 299260 50396 299266
rect 50344 299202 50396 299208
rect 43444 299124 43496 299130
rect 43444 299066 43496 299072
rect 40684 255264 40736 255270
rect 40684 255206 40736 255212
rect 39396 241460 39448 241466
rect 39396 241402 39448 241408
rect 39304 85536 39356 85542
rect 39304 85478 39356 85484
rect 39304 39364 39356 39370
rect 39304 39306 39356 39312
rect 37188 7608 37240 7614
rect 37188 7550 37240 7556
rect 35164 4072 35216 4078
rect 35164 4014 35216 4020
rect 34796 4004 34848 4010
rect 34796 3946 34848 3952
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 34808 480 34836 3946
rect 35992 3868 36044 3874
rect 35992 3810 36044 3816
rect 36004 480 36032 3810
rect 37200 480 37228 7550
rect 38384 4072 38436 4078
rect 38384 4014 38436 4020
rect 38396 480 38424 4014
rect 39316 3942 39344 39306
rect 40684 7676 40736 7682
rect 40684 7618 40736 7624
rect 39304 3936 39356 3942
rect 39304 3878 39356 3884
rect 39580 3392 39632 3398
rect 39580 3334 39632 3340
rect 39592 480 39620 3334
rect 40696 480 40724 7618
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 41880 3324 41932 3330
rect 41880 3266 41932 3272
rect 41892 480 41920 3266
rect 43088 480 43116 3878
rect 43456 3398 43484 299066
rect 47584 296064 47636 296070
rect 47584 296006 47636 296012
rect 44272 7744 44324 7750
rect 44272 7686 44324 7692
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 44284 480 44312 7686
rect 47596 4078 47624 296006
rect 48964 7812 49016 7818
rect 48964 7754 49016 7760
rect 47860 5500 47912 5506
rect 47860 5442 47912 5448
rect 47584 4072 47636 4078
rect 47584 4014 47636 4020
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45480 480 45508 3334
rect 46664 3052 46716 3058
rect 46664 2994 46716 3000
rect 46676 480 46704 2994
rect 47872 480 47900 5442
rect 48976 480 49004 7754
rect 50160 3324 50212 3330
rect 50160 3266 50212 3272
rect 50172 480 50200 3266
rect 50356 3058 50384 299202
rect 51736 293962 51764 701791
rect 61384 700596 61436 700602
rect 61384 700538 61436 700544
rect 57244 297492 57296 297498
rect 57244 297434 57296 297440
rect 54484 296132 54536 296138
rect 54484 296074 54536 296080
rect 51816 294704 51868 294710
rect 51816 294646 51868 294652
rect 51724 293956 51776 293962
rect 51724 293898 51776 293904
rect 51356 4752 51408 4758
rect 51356 4694 51408 4700
rect 50344 3052 50396 3058
rect 50344 2994 50396 3000
rect 51368 480 51396 4694
rect 51828 4010 51856 294646
rect 52552 7880 52604 7886
rect 52552 7822 52604 7828
rect 51816 4004 51868 4010
rect 51816 3946 51868 3952
rect 52564 480 52592 7822
rect 53748 4004 53800 4010
rect 53748 3946 53800 3952
rect 53760 480 53788 3946
rect 54496 3398 54524 296074
rect 56048 7948 56100 7954
rect 56048 7890 56100 7896
rect 54944 4684 54996 4690
rect 54944 4626 54996 4632
rect 54484 3392 54536 3398
rect 54484 3334 54536 3340
rect 54956 480 54984 4626
rect 56060 480 56088 7890
rect 57256 4078 57284 297434
rect 61396 45558 61424 700538
rect 72988 700262 73016 703520
rect 89180 700330 89208 703520
rect 105464 700777 105492 703520
rect 137284 701412 137336 701418
rect 137284 701354 137336 701360
rect 105450 700768 105506 700777
rect 105450 700703 105506 700712
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 72976 700256 73028 700262
rect 72976 700198 73028 700204
rect 107568 299464 107620 299470
rect 107568 299406 107620 299412
rect 103428 299396 103480 299402
rect 103428 299338 103480 299344
rect 90364 299328 90416 299334
rect 90364 299270 90416 299276
rect 87604 298512 87656 298518
rect 87604 298454 87656 298460
rect 83464 298444 83516 298450
rect 83464 298386 83516 298392
rect 79324 298376 79376 298382
rect 79324 298318 79376 298324
rect 61384 45552 61436 45558
rect 61384 45494 61436 45500
rect 73804 8288 73856 8294
rect 73804 8230 73856 8236
rect 70308 8220 70360 8226
rect 70308 8162 70360 8168
rect 66720 8152 66772 8158
rect 66720 8094 66772 8100
rect 63224 8084 63276 8090
rect 63224 8026 63276 8032
rect 59636 8016 59688 8022
rect 59636 7958 59688 7964
rect 58440 4548 58492 4554
rect 58440 4490 58492 4496
rect 57244 4072 57296 4078
rect 57244 4014 57296 4020
rect 57244 3256 57296 3262
rect 57244 3198 57296 3204
rect 57256 480 57284 3198
rect 58452 480 58480 4490
rect 59648 480 59676 7958
rect 62028 4616 62080 4622
rect 62028 4558 62080 4564
rect 60832 4072 60884 4078
rect 60832 4014 60884 4020
rect 60844 480 60872 4014
rect 62040 480 62068 4558
rect 63236 480 63264 8026
rect 65524 4480 65576 4486
rect 65524 4422 65576 4428
rect 64328 3188 64380 3194
rect 64328 3130 64380 3136
rect 64340 480 64368 3130
rect 65536 480 65564 4422
rect 66732 480 66760 8094
rect 69112 4344 69164 4350
rect 69112 4286 69164 4292
rect 67916 4140 67968 4146
rect 67916 4082 67968 4088
rect 67928 480 67956 4082
rect 69124 480 69152 4286
rect 70320 480 70348 8162
rect 72608 4412 72660 4418
rect 72608 4354 72660 4360
rect 71504 3120 71556 3126
rect 71504 3062 71556 3068
rect 71516 480 71544 3062
rect 72620 480 72648 4354
rect 73816 480 73844 8230
rect 77392 7540 77444 7546
rect 77392 7482 77444 7488
rect 76196 4276 76248 4282
rect 76196 4218 76248 4224
rect 75000 3392 75052 3398
rect 75000 3334 75052 3340
rect 75012 480 75040 3334
rect 76208 480 76236 4218
rect 77404 480 77432 7482
rect 79336 3330 79364 298318
rect 81348 14476 81400 14482
rect 81348 14418 81400 14424
rect 79692 6316 79744 6322
rect 79692 6258 79744 6264
rect 79324 3324 79376 3330
rect 79324 3266 79376 3272
rect 78588 3052 78640 3058
rect 78588 2994 78640 3000
rect 78600 480 78628 2994
rect 79704 480 79732 6258
rect 81360 3330 81388 14418
rect 83280 6384 83332 6390
rect 83280 6326 83332 6332
rect 80888 3324 80940 3330
rect 80888 3266 80940 3272
rect 81348 3324 81400 3330
rect 81348 3266 81400 3272
rect 80900 480 80928 3266
rect 82084 2984 82136 2990
rect 82084 2926 82136 2932
rect 82096 480 82124 2926
rect 83292 480 83320 6326
rect 83476 3262 83504 298386
rect 86224 297560 86276 297566
rect 86224 297502 86276 297508
rect 86236 3330 86264 297502
rect 86868 6452 86920 6458
rect 86868 6394 86920 6400
rect 84476 3324 84528 3330
rect 84476 3266 84528 3272
rect 86224 3324 86276 3330
rect 86224 3266 86276 3272
rect 83464 3256 83516 3262
rect 83464 3198 83516 3204
rect 84488 480 84516 3266
rect 85672 3256 85724 3262
rect 85672 3198 85724 3204
rect 85684 480 85712 3198
rect 86880 480 86908 6394
rect 87616 3194 87644 298454
rect 88984 297628 89036 297634
rect 88984 297570 89036 297576
rect 88996 3330 89024 297570
rect 90376 3330 90404 299270
rect 101404 298716 101456 298722
rect 101404 298658 101456 298664
rect 98644 298308 98696 298314
rect 98644 298250 98696 298256
rect 93124 297696 93176 297702
rect 93124 297638 93176 297644
rect 90456 6520 90508 6526
rect 90456 6462 90508 6468
rect 87972 3324 88024 3330
rect 87972 3266 88024 3272
rect 88984 3324 89036 3330
rect 88984 3266 89036 3272
rect 89168 3324 89220 3330
rect 89168 3266 89220 3272
rect 90364 3324 90416 3330
rect 90364 3266 90416 3272
rect 87604 3188 87656 3194
rect 87604 3130 87656 3136
rect 87984 480 88012 3266
rect 89180 480 89208 3266
rect 90468 3210 90496 6462
rect 93136 3330 93164 297638
rect 95148 296200 95200 296206
rect 95148 296142 95200 296148
rect 93952 6588 94004 6594
rect 93952 6530 94004 6536
rect 91560 3324 91612 3330
rect 91560 3266 91612 3272
rect 93124 3324 93176 3330
rect 93124 3266 93176 3272
rect 90376 3182 90496 3210
rect 90376 480 90404 3182
rect 91572 480 91600 3266
rect 92756 3188 92808 3194
rect 92756 3130 92808 3136
rect 92768 480 92796 3130
rect 93964 480 93992 6530
rect 95160 480 95188 296142
rect 98656 6914 98684 298250
rect 99288 296268 99340 296274
rect 99288 296210 99340 296216
rect 98564 6886 98684 6914
rect 97448 6656 97500 6662
rect 97448 6598 97500 6604
rect 96252 2984 96304 2990
rect 96252 2926 96304 2932
rect 96264 480 96292 2926
rect 97460 480 97488 6598
rect 98564 3126 98592 6886
rect 99300 3126 99328 296210
rect 101036 7472 101088 7478
rect 101036 7414 101088 7420
rect 98552 3120 98604 3126
rect 98552 3062 98604 3068
rect 98644 3120 98696 3126
rect 98644 3062 98696 3068
rect 99288 3120 99340 3126
rect 99288 3062 99340 3068
rect 98656 480 98684 3062
rect 99840 3052 99892 3058
rect 99840 2994 99892 3000
rect 99852 480 99880 2994
rect 101048 480 101076 7414
rect 101416 2990 101444 298658
rect 103440 6914 103468 299338
rect 105544 298240 105596 298246
rect 105544 298182 105596 298188
rect 104164 297764 104216 297770
rect 104164 297706 104216 297712
rect 103348 6886 103468 6914
rect 102232 3120 102284 3126
rect 102232 3062 102284 3068
rect 101404 2984 101456 2990
rect 101404 2926 101456 2932
rect 102244 480 102272 3062
rect 103348 480 103376 6886
rect 104176 3126 104204 297706
rect 104532 8968 104584 8974
rect 104532 8910 104584 8916
rect 104164 3120 104216 3126
rect 104164 3062 104216 3068
rect 104544 480 104572 8910
rect 105556 2922 105584 298182
rect 107580 3126 107608 299406
rect 114468 298648 114520 298654
rect 114468 298590 114520 298596
rect 111064 297832 111116 297838
rect 111064 297774 111116 297780
rect 108304 296336 108356 296342
rect 108304 296278 108356 296284
rect 108120 9104 108172 9110
rect 108120 9046 108172 9052
rect 106924 3120 106976 3126
rect 106924 3062 106976 3068
rect 107568 3120 107620 3126
rect 107568 3062 107620 3068
rect 105728 2984 105780 2990
rect 105728 2926 105780 2932
rect 105544 2916 105596 2922
rect 105544 2858 105596 2864
rect 105740 480 105768 2926
rect 106936 480 106964 3062
rect 108132 480 108160 9046
rect 108316 2990 108344 296278
rect 111076 3126 111104 297774
rect 113088 296404 113140 296410
rect 113088 296346 113140 296352
rect 111616 9036 111668 9042
rect 111616 8978 111668 8984
rect 109316 3120 109368 3126
rect 109316 3062 109368 3068
rect 111064 3120 111116 3126
rect 111064 3062 111116 3068
rect 108304 2984 108356 2990
rect 108304 2926 108356 2932
rect 109328 480 109356 3062
rect 110512 2984 110564 2990
rect 110512 2926 110564 2932
rect 110524 480 110552 2926
rect 111628 480 111656 8978
rect 113100 6914 113128 296346
rect 112824 6886 113128 6914
rect 112824 480 112852 6886
rect 114480 2990 114508 298590
rect 121368 298580 121420 298586
rect 121368 298522 121420 298528
rect 117228 294840 117280 294846
rect 117228 294782 117280 294788
rect 115204 9172 115256 9178
rect 115204 9114 115256 9120
rect 114008 2984 114060 2990
rect 114008 2926 114060 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 114020 480 114048 2926
rect 115216 480 115244 9114
rect 117240 2990 117268 294782
rect 119988 294772 120040 294778
rect 119988 294714 120040 294720
rect 119804 10396 119856 10402
rect 119804 10338 119856 10344
rect 119816 2990 119844 10338
rect 120000 6914 120028 294714
rect 121380 6914 121408 298522
rect 135168 298036 135220 298042
rect 135168 297978 135220 297984
rect 133788 297968 133840 297974
rect 133788 297910 133840 297916
rect 129648 297900 129700 297906
rect 129648 297842 129700 297848
rect 124128 294908 124180 294914
rect 124128 294850 124180 294856
rect 122748 10464 122800 10470
rect 122748 10406 122800 10412
rect 119908 6886 120028 6914
rect 121104 6886 121408 6914
rect 116400 2984 116452 2990
rect 116400 2926 116452 2932
rect 117228 2984 117280 2990
rect 117228 2926 117280 2932
rect 118792 2984 118844 2990
rect 118792 2926 118844 2932
rect 119804 2984 119856 2990
rect 119804 2926 119856 2932
rect 116412 480 116440 2926
rect 117596 2916 117648 2922
rect 117596 2858 117648 2864
rect 117608 480 117636 2858
rect 118804 480 118832 2926
rect 119908 480 119936 6886
rect 121104 480 121132 6886
rect 122760 2990 122788 10406
rect 124140 2990 124168 294850
rect 126888 10600 126940 10606
rect 126888 10542 126940 10548
rect 126900 2990 126928 10542
rect 128176 7404 128228 7410
rect 128176 7346 128228 7352
rect 126980 6724 127032 6730
rect 126980 6666 127032 6672
rect 122288 2984 122340 2990
rect 122288 2926 122340 2932
rect 122748 2984 122800 2990
rect 122748 2926 122800 2932
rect 123484 2984 123536 2990
rect 123484 2926 123536 2932
rect 124128 2984 124180 2990
rect 124128 2926 124180 2932
rect 125876 2984 125928 2990
rect 125876 2926 125928 2932
rect 126888 2984 126940 2990
rect 126888 2926 126940 2932
rect 122300 480 122328 2926
rect 123496 480 123524 2926
rect 124680 2848 124732 2854
rect 124680 2790 124732 2796
rect 124692 480 124720 2790
rect 125888 480 125916 2926
rect 126992 480 127020 6666
rect 128188 480 128216 7346
rect 129660 6914 129688 297842
rect 132408 12028 132460 12034
rect 132408 11970 132460 11976
rect 129384 6886 129688 6914
rect 129384 480 129412 6886
rect 130568 6792 130620 6798
rect 130568 6734 130620 6740
rect 130580 480 130608 6734
rect 132420 2854 132448 11970
rect 133800 2854 133828 297910
rect 135180 2854 135208 297978
rect 137296 202842 137324 701354
rect 137848 701010 137876 703520
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 154132 700913 154160 703520
rect 154118 700904 154174 700913
rect 154118 700839 154174 700848
rect 170324 700641 170352 703520
rect 182180 703452 182232 703458
rect 182180 703394 182232 703400
rect 180064 702704 180116 702710
rect 180064 702646 180116 702652
rect 170310 700632 170366 700641
rect 170310 700567 170366 700576
rect 177302 700224 177358 700233
rect 177302 700159 177358 700168
rect 177316 346390 177344 700159
rect 177304 346384 177356 346390
rect 177304 346326 177356 346332
rect 140688 298104 140740 298110
rect 140688 298046 140740 298052
rect 137284 202836 137336 202842
rect 137284 202778 137336 202784
rect 137928 202156 137980 202162
rect 137928 202098 137980 202104
rect 136456 10532 136508 10538
rect 136456 10474 136508 10480
rect 135260 9240 135312 9246
rect 135260 9182 135312 9188
rect 131764 2848 131816 2854
rect 131764 2790 131816 2796
rect 132408 2848 132460 2854
rect 132408 2790 132460 2796
rect 132960 2848 133012 2854
rect 132960 2790 133012 2796
rect 133788 2848 133840 2854
rect 133788 2790 133840 2796
rect 134156 2848 134208 2854
rect 134156 2790 134208 2796
rect 135168 2848 135220 2854
rect 135168 2790 135220 2796
rect 131776 480 131804 2790
rect 132972 480 133000 2790
rect 134168 480 134196 2790
rect 135272 480 135300 9182
rect 136468 480 136496 10474
rect 137940 6914 137968 202098
rect 138848 9308 138900 9314
rect 138848 9250 138900 9256
rect 137664 6886 137968 6914
rect 137664 480 137692 6886
rect 138860 480 138888 9250
rect 140700 2854 140728 298046
rect 179328 297356 179380 297362
rect 179328 297298 179380 297304
rect 144828 297288 144880 297294
rect 144828 297230 144880 297236
rect 142068 297220 142120 297226
rect 142068 297162 142120 297168
rect 142080 2854 142108 297162
rect 144736 11756 144788 11762
rect 144736 11698 144788 11704
rect 142436 9376 142488 9382
rect 142436 9318 142488 9324
rect 140044 2848 140096 2854
rect 140044 2790 140096 2796
rect 140688 2848 140740 2854
rect 140688 2790 140740 2796
rect 141240 2848 141292 2854
rect 141240 2790 141292 2796
rect 142068 2848 142120 2854
rect 142068 2790 142120 2796
rect 140056 480 140084 2790
rect 141252 480 141280 2790
rect 142448 480 142476 9318
rect 143540 2848 143592 2854
rect 143540 2790 143592 2796
rect 143552 480 143580 2790
rect 144748 480 144776 11698
rect 144840 2854 144868 297230
rect 177948 296676 178000 296682
rect 177948 296618 178000 296624
rect 158628 296608 158680 296614
rect 158628 296550 158680 296556
rect 147588 296540 147640 296546
rect 147588 296482 147640 296488
rect 145932 9444 145984 9450
rect 145932 9386 145984 9392
rect 144828 2848 144880 2854
rect 144828 2790 144880 2796
rect 145944 480 145972 9386
rect 147600 2854 147628 296482
rect 151728 296472 151780 296478
rect 151728 296414 151780 296420
rect 148968 295928 149020 295934
rect 148968 295870 149020 295876
rect 148980 2854 149008 295870
rect 149520 9580 149572 9586
rect 149520 9522 149572 9528
rect 147128 2848 147180 2854
rect 147128 2790 147180 2796
rect 147588 2848 147640 2854
rect 147588 2790 147640 2796
rect 148324 2848 148376 2854
rect 148324 2790 148376 2796
rect 148968 2848 149020 2854
rect 148968 2790 149020 2796
rect 147140 480 147168 2790
rect 148336 480 148364 2790
rect 149532 480 149560 9522
rect 151740 2854 151768 296414
rect 153108 188352 153160 188358
rect 153108 188294 153160 188300
rect 153016 9512 153068 9518
rect 153016 9454 153068 9460
rect 150624 2848 150676 2854
rect 150624 2790 150676 2796
rect 151728 2848 151780 2854
rect 151728 2790 151780 2796
rect 151820 2848 151872 2854
rect 151820 2790 151872 2796
rect 150636 480 150664 2790
rect 151832 480 151860 2790
rect 153028 480 153056 9454
rect 153120 2854 153148 188294
rect 155868 49020 155920 49026
rect 155868 48962 155920 48968
rect 154212 11824 154264 11830
rect 154212 11766 154264 11772
rect 153108 2848 153160 2854
rect 153108 2790 153160 2796
rect 154224 480 154252 11766
rect 155880 2854 155908 48962
rect 156604 9648 156656 9654
rect 156604 9590 156656 9596
rect 155408 2848 155460 2854
rect 155408 2790 155460 2796
rect 155868 2848 155920 2854
rect 155868 2790 155920 2796
rect 155420 480 155448 2790
rect 156616 480 156644 9590
rect 158640 2854 158668 296550
rect 169668 13184 169720 13190
rect 169668 13126 169720 13132
rect 161296 10940 161348 10946
rect 161296 10882 161348 10888
rect 160100 8900 160152 8906
rect 160100 8842 160152 8848
rect 158904 7336 158956 7342
rect 158904 7278 158956 7284
rect 157800 2848 157852 2854
rect 157800 2790 157852 2796
rect 158628 2848 158680 2854
rect 158628 2790 158680 2796
rect 157812 480 157840 2790
rect 158916 480 158944 7278
rect 160112 480 160140 8842
rect 161308 480 161336 10882
rect 165528 10872 165580 10878
rect 165528 10814 165580 10820
rect 163688 7268 163740 7274
rect 163688 7210 163740 7216
rect 162492 6860 162544 6866
rect 162492 6802 162544 6808
rect 162504 480 162532 6802
rect 163700 480 163728 7210
rect 165540 2854 165568 10814
rect 167184 7200 167236 7206
rect 167184 7142 167236 7148
rect 166080 6112 166132 6118
rect 166080 6054 166132 6060
rect 164884 2848 164936 2854
rect 164884 2790 164936 2796
rect 165528 2848 165580 2854
rect 165528 2790 165580 2796
rect 164896 480 164924 2790
rect 166092 480 166120 6054
rect 167196 480 167224 7142
rect 169576 6044 169628 6050
rect 169576 5986 169628 5992
rect 168380 2848 168432 2854
rect 168380 2790 168432 2796
rect 168392 480 168420 2790
rect 169588 480 169616 5986
rect 169680 2854 169708 13126
rect 176568 11892 176620 11898
rect 176568 11834 176620 11840
rect 172428 10260 172480 10266
rect 172428 10202 172480 10208
rect 170772 7132 170824 7138
rect 170772 7074 170824 7080
rect 169668 2848 169720 2854
rect 169668 2790 169720 2796
rect 170784 480 170812 7074
rect 172440 2854 172468 10202
rect 174268 7064 174320 7070
rect 174268 7006 174320 7012
rect 173164 5976 173216 5982
rect 173164 5918 173216 5924
rect 171968 2848 172020 2854
rect 171968 2790 172020 2796
rect 172428 2848 172480 2854
rect 172428 2790 172480 2796
rect 171980 480 172008 2790
rect 173176 480 173204 5918
rect 174280 480 174308 7006
rect 176580 2854 176608 11834
rect 177960 6914 177988 296618
rect 179340 6914 179368 297298
rect 180076 164218 180104 702646
rect 181812 701752 181864 701758
rect 181812 701694 181864 701700
rect 181824 302938 181852 701694
rect 182088 701684 182140 701690
rect 182088 701626 182140 701632
rect 181904 701616 181956 701622
rect 181904 701558 181956 701564
rect 181812 302932 181864 302938
rect 181812 302874 181864 302880
rect 180064 164212 180116 164218
rect 180064 164154 180116 164160
rect 181916 73166 181944 701558
rect 181996 701140 182048 701146
rect 181996 701082 182048 701088
rect 181904 73160 181956 73166
rect 181904 73102 181956 73108
rect 182008 33114 182036 701082
rect 181996 33108 182048 33114
rect 181996 33050 182048 33056
rect 182100 20602 182128 701626
rect 182192 684486 182220 703394
rect 182272 703316 182324 703322
rect 182272 703258 182324 703264
rect 182180 684480 182232 684486
rect 182180 684422 182232 684428
rect 182284 633418 182312 703258
rect 182364 703248 182416 703254
rect 182364 703190 182416 703196
rect 182272 633412 182324 633418
rect 182272 633354 182324 633360
rect 182376 580990 182404 703190
rect 182456 703180 182508 703186
rect 182456 703122 182508 703128
rect 182364 580984 182416 580990
rect 182364 580926 182416 580932
rect 182468 528562 182496 703122
rect 182548 703112 182600 703118
rect 182548 703054 182600 703060
rect 182456 528556 182508 528562
rect 182456 528498 182508 528504
rect 182560 476066 182588 703054
rect 182640 703044 182692 703050
rect 182640 702986 182692 702992
rect 182548 476060 182600 476066
rect 182548 476002 182600 476008
rect 182652 423638 182680 702986
rect 182732 702976 182784 702982
rect 182732 702918 182784 702924
rect 182640 423632 182692 423638
rect 182640 423574 182692 423580
rect 182744 372570 182772 702918
rect 201696 701690 202078 701706
rect 201684 701684 202078 701690
rect 201736 701678 202078 701684
rect 201684 701626 201736 701632
rect 191196 701616 191248 701622
rect 191248 701564 191590 701570
rect 191196 701558 191590 701564
rect 183008 701548 183060 701554
rect 191208 701542 191590 701558
rect 183008 701490 183060 701496
rect 182916 701480 182968 701486
rect 182916 701422 182968 701428
rect 182824 701072 182876 701078
rect 182824 701014 182876 701020
rect 182732 372564 182784 372570
rect 182732 372506 182784 372512
rect 182732 318844 182784 318850
rect 182732 318786 182784 318792
rect 182744 303521 182772 318786
rect 182730 303512 182786 303521
rect 182730 303447 182786 303456
rect 182836 303006 182864 701014
rect 182824 303000 182876 303006
rect 182824 302942 182876 302948
rect 182180 299532 182232 299538
rect 182180 299474 182232 299480
rect 182088 20596 182140 20602
rect 182088 20538 182140 20544
rect 182088 11960 182140 11966
rect 182088 11902 182140 11908
rect 177868 6886 177988 6914
rect 179064 6886 179368 6914
rect 176660 5908 176712 5914
rect 176660 5850 176712 5856
rect 175464 2848 175516 2854
rect 175464 2790 175516 2796
rect 176568 2848 176620 2854
rect 176568 2790 176620 2796
rect 175476 480 175504 2790
rect 176672 480 176700 5850
rect 177868 480 177896 6886
rect 179064 480 179092 6886
rect 180248 5840 180300 5846
rect 180248 5782 180300 5788
rect 180260 480 180288 5782
rect 182100 3534 182128 11902
rect 182192 4894 182220 299474
rect 182928 113150 182956 701422
rect 182916 113144 182968 113150
rect 182916 113086 182968 113092
rect 183020 86970 183048 701490
rect 183100 701208 183152 701214
rect 194692 701208 194744 701214
rect 183100 701150 183152 701156
rect 183008 86964 183060 86970
rect 183008 86906 183060 86912
rect 183112 46918 183140 701150
rect 184216 701134 184598 701162
rect 187712 701146 188094 701162
rect 194744 701156 195086 701162
rect 194692 701150 195086 701156
rect 187700 701140 188094 701146
rect 184216 701078 184244 701134
rect 187752 701134 188094 701140
rect 194704 701134 195086 701150
rect 198200 701146 198582 701162
rect 198188 701140 198582 701146
rect 187700 701082 187752 701088
rect 198240 701134 198582 701140
rect 198188 701082 198240 701088
rect 202800 701078 202828 703520
rect 218992 702001 219020 703520
rect 235184 703474 235212 703520
rect 235368 703474 235396 703582
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 310886 703624 310942 703633
rect 300308 703588 300360 703594
rect 310886 703559 310942 703568
rect 300308 703530 300360 703536
rect 235184 703446 235396 703474
rect 258172 702908 258224 702914
rect 258172 702850 258224 702856
rect 254676 702840 254728 702846
rect 254676 702782 254728 702788
rect 226616 702772 226668 702778
rect 226616 702714 226668 702720
rect 219624 702636 219676 702642
rect 219624 702578 219676 702584
rect 212630 701992 212686 702001
rect 212630 701927 212686 701936
rect 216126 701992 216182 702001
rect 216126 701927 216182 701936
rect 218978 701992 219034 702001
rect 218978 701927 219034 701936
rect 212644 701692 212672 701927
rect 216140 701692 216168 701927
rect 219636 701692 219664 702578
rect 223118 701992 223174 702001
rect 223118 701927 223174 701936
rect 223132 701692 223160 701927
rect 226628 701692 226656 702714
rect 251178 702536 251234 702545
rect 251178 702471 251234 702480
rect 244002 702400 244058 702409
rect 244002 702335 244058 702344
rect 247682 702400 247738 702409
rect 247682 702335 247738 702344
rect 247866 702400 247922 702409
rect 247866 702335 247922 702344
rect 233606 702128 233662 702137
rect 233606 702063 233662 702072
rect 240690 702128 240746 702137
rect 240690 702063 240746 702072
rect 230110 701992 230166 702001
rect 230110 701927 230166 701936
rect 230124 701692 230152 701927
rect 233620 701692 233648 702063
rect 237194 701992 237250 702001
rect 237194 701927 237250 701936
rect 237208 701692 237236 701927
rect 240704 701692 240732 702063
rect 205192 701554 205574 701570
rect 205180 701548 205574 701554
rect 205232 701542 205574 701548
rect 205180 701490 205232 701496
rect 208676 701480 208728 701486
rect 208728 701428 209070 701434
rect 208676 701422 209070 701428
rect 208688 701406 209070 701422
rect 244016 701418 244044 702335
rect 244186 702264 244242 702273
rect 244186 702199 244242 702208
rect 244200 701692 244228 702199
rect 247696 701692 247724 702335
rect 244004 701412 244056 701418
rect 244004 701354 244056 701360
rect 247880 701350 247908 702335
rect 251192 701692 251220 702471
rect 254688 701692 254716 702782
rect 258184 701692 258212 702850
rect 247868 701344 247920 701350
rect 247868 701286 247920 701292
rect 261786 701134 262076 701162
rect 265282 701134 265664 701162
rect 262048 701078 262076 701134
rect 265636 701078 265664 701134
rect 267660 701078 267688 703520
rect 268752 702092 268804 702098
rect 268752 702034 268804 702040
rect 268764 701692 268792 702034
rect 282762 701554 282868 701570
rect 282762 701548 282880 701554
rect 282762 701542 282828 701548
rect 282828 701490 282880 701496
rect 279608 701480 279660 701486
rect 275770 701418 275968 701434
rect 279266 701428 279608 701434
rect 279266 701422 279660 701428
rect 275770 701412 275980 701418
rect 275770 701406 275928 701412
rect 279266 701406 279648 701422
rect 275928 701354 275980 701360
rect 272616 701344 272668 701350
rect 272274 701292 272616 701298
rect 272274 701286 272668 701292
rect 272274 701270 272656 701286
rect 283852 701078 283880 703520
rect 300136 703474 300164 703520
rect 300320 703474 300348 703530
rect 300136 703446 300348 703474
rect 300308 702568 300360 702574
rect 300308 702510 300360 702516
rect 289820 702228 289872 702234
rect 289820 702170 289872 702176
rect 289832 701692 289860 702170
rect 297088 701752 297140 701758
rect 293342 701690 293632 701706
rect 296838 701700 297088 701706
rect 296838 701694 297140 701700
rect 293342 701684 293644 701690
rect 293342 701678 293592 701684
rect 296838 701678 297128 701694
rect 300320 701692 300348 702510
rect 307300 701888 307352 701894
rect 307300 701830 307352 701836
rect 304080 701820 304132 701826
rect 304080 701762 304132 701768
rect 304092 701706 304120 701762
rect 303830 701678 304120 701706
rect 307312 701692 307340 701830
rect 310900 701692 310928 703559
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 363512 703656 363564 703662
rect 363512 703598 363564 703604
rect 321374 703488 321430 703497
rect 321374 703423 321430 703432
rect 316130 702536 316186 702545
rect 316130 702471 316186 702480
rect 314384 702160 314436 702166
rect 314384 702102 314436 702108
rect 314396 701692 314424 702102
rect 293592 701626 293644 701632
rect 286600 701616 286652 701622
rect 286350 701564 286600 701570
rect 286350 701558 286652 701564
rect 286350 701542 286640 701558
rect 316144 701146 316172 702471
rect 321388 701692 321416 703423
rect 331862 702944 331918 702953
rect 331862 702879 331918 702888
rect 328368 702024 328420 702030
rect 328368 701966 328420 701972
rect 324872 701956 324924 701962
rect 324872 701898 324924 701904
rect 324884 701692 324912 701898
rect 328380 701692 328408 701966
rect 331876 701692 331904 702879
rect 316132 701140 316184 701146
rect 317906 701134 318288 701162
rect 316132 701082 316184 701088
rect 318260 701078 318288 701134
rect 332520 701078 332548 703520
rect 348804 703474 348832 703520
rect 348974 703488 349030 703497
rect 348804 703446 348974 703474
rect 348974 703423 349030 703432
rect 353298 703488 353354 703497
rect 353298 703423 353354 703432
rect 349436 703384 349488 703390
rect 349436 703326 349488 703332
rect 342442 702808 342498 702817
rect 342442 702743 342498 702752
rect 333978 702672 334034 702681
rect 333978 702607 334034 702616
rect 333242 702536 333298 702545
rect 333242 702471 333298 702480
rect 333256 701078 333284 702471
rect 333992 702234 334020 702607
rect 333980 702228 334032 702234
rect 333980 702170 334032 702176
rect 338948 702228 339000 702234
rect 338948 702170 339000 702176
rect 338960 701692 338988 702170
rect 342456 701692 342484 702743
rect 345938 702536 345994 702545
rect 345938 702471 345994 702480
rect 349066 702536 349122 702545
rect 349066 702471 349122 702480
rect 345952 701692 345980 702471
rect 335478 701146 335768 701162
rect 335478 701140 335780 701146
rect 335478 701134 335728 701140
rect 335728 701082 335780 701088
rect 349080 701078 349108 702471
rect 349448 701692 349476 703326
rect 353312 702817 353340 703423
rect 362958 703080 363014 703089
rect 362958 703015 363014 703024
rect 353114 702808 353170 702817
rect 353114 702743 353170 702752
rect 353298 702808 353354 702817
rect 353298 702743 353354 702752
rect 353128 702545 353156 702743
rect 362222 702672 362278 702681
rect 362222 702607 362278 702616
rect 352930 702536 352986 702545
rect 352930 702471 352986 702480
rect 353114 702536 353170 702545
rect 353114 702471 353170 702480
rect 352944 701692 352972 702471
rect 362236 701214 362264 702607
rect 362972 701214 363000 703015
rect 363524 701692 363552 703598
rect 364954 703520 365066 704960
rect 365718 703896 365774 703905
rect 365718 703831 365774 703840
rect 374642 703896 374698 703905
rect 374642 703831 374698 703840
rect 364996 701214 365024 703520
rect 365732 702506 365760 703831
rect 374552 703520 374604 703526
rect 374552 703462 374604 703468
rect 369674 703080 369730 703089
rect 369674 703015 369730 703024
rect 369688 702681 369716 703015
rect 369490 702672 369546 702681
rect 369490 702607 369546 702616
rect 369674 702672 369730 702681
rect 369674 702607 369730 702616
rect 365810 702536 365866 702545
rect 365720 702500 365772 702506
rect 365810 702471 365866 702480
rect 365720 702442 365772 702448
rect 362224 701208 362276 701214
rect 356454 701134 356744 701162
rect 360042 701134 360148 701162
rect 362224 701150 362276 701156
rect 362960 701208 363012 701214
rect 362960 701150 363012 701156
rect 364984 701208 365036 701214
rect 364984 701150 365036 701156
rect 365824 701146 365852 702471
rect 367100 701208 367152 701214
rect 367034 701156 367100 701162
rect 367034 701150 367152 701156
rect 356716 701078 356744 701134
rect 360120 701078 360148 701134
rect 365812 701140 365864 701146
rect 367034 701134 367140 701150
rect 369504 701146 369532 702607
rect 369674 702536 369730 702545
rect 374090 702536 374146 702545
rect 369674 702471 369676 702480
rect 369728 702471 369730 702480
rect 370504 702500 370556 702506
rect 369676 702442 369728 702448
rect 374090 702471 374146 702480
rect 370504 702442 370556 702448
rect 370516 701692 370544 702442
rect 373828 701146 374026 701162
rect 374104 701146 374132 702471
rect 374564 702098 374592 703462
rect 374656 703089 374684 703831
rect 381146 703520 381258 704960
rect 395066 703760 395122 703769
rect 395066 703695 395122 703704
rect 384580 703588 384632 703594
rect 384580 703530 384632 703536
rect 374642 703080 374698 703089
rect 374642 703015 374698 703024
rect 375380 702568 375432 702574
rect 375380 702510 375432 702516
rect 380990 702536 381046 702545
rect 375392 702409 375420 702510
rect 380990 702471 381046 702480
rect 374642 702400 374698 702409
rect 374642 702335 374698 702344
rect 375378 702400 375434 702409
rect 375378 702335 375434 702344
rect 374656 702098 374684 702335
rect 374552 702092 374604 702098
rect 374552 702034 374604 702040
rect 374644 702092 374696 702098
rect 374644 702034 374696 702040
rect 381004 701692 381032 702471
rect 384592 701692 384620 703530
rect 391110 702536 391166 702545
rect 391110 702471 391166 702480
rect 391124 701214 391152 702471
rect 395080 701692 395108 703695
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429660 703656 429712 703662
rect 429660 703598 429712 703604
rect 391112 701208 391164 701214
rect 377232 701146 377522 701162
rect 387812 701146 388102 701162
rect 391112 701150 391164 701156
rect 391216 701146 391598 701162
rect 397472 701146 397500 703520
rect 405554 703488 405610 703497
rect 405554 703423 405610 703432
rect 404360 702568 404412 702574
rect 404360 702510 404412 702516
rect 369492 701140 369544 701146
rect 365812 701082 365864 701088
rect 369492 701082 369544 701088
rect 373816 701140 374026 701146
rect 373868 701134 374026 701140
rect 374092 701140 374144 701146
rect 373816 701082 373868 701088
rect 374092 701082 374144 701088
rect 377220 701140 377522 701146
rect 377272 701134 377522 701140
rect 387800 701140 388102 701146
rect 377220 701082 377272 701088
rect 387852 701134 388102 701140
rect 391204 701140 391598 701146
rect 387800 701082 387852 701088
rect 391256 701134 391598 701140
rect 397460 701140 397512 701146
rect 391204 701082 391256 701088
rect 397460 701082 397512 701088
rect 398208 701134 398590 701162
rect 401704 701134 402086 701162
rect 398208 701078 398236 701134
rect 401704 701078 401732 701134
rect 404372 701078 404400 702510
rect 405568 701692 405596 703423
rect 412638 702672 412694 702681
rect 412638 702607 412694 702616
rect 409052 702568 409104 702574
rect 409052 702510 409104 702516
rect 409064 701692 409092 702510
rect 412652 701692 412680 702607
rect 413664 702506 413692 703520
rect 429672 703474 429700 703598
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 552940 703792 552992 703798
rect 552940 703734 552992 703740
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 437204 703452 437256 703458
rect 437204 703394 437256 703400
rect 426622 703352 426678 703361
rect 426622 703287 426678 703296
rect 416134 703216 416190 703225
rect 416134 703151 416190 703160
rect 418066 703216 418122 703225
rect 418066 703151 418122 703160
rect 413652 702500 413704 702506
rect 413652 702442 413704 702448
rect 416148 701692 416176 703151
rect 418080 702166 418108 703151
rect 418068 702160 418120 702166
rect 418068 702102 418120 702108
rect 426636 701692 426664 703287
rect 427634 702672 427690 702681
rect 427634 702607 427690 702616
rect 427648 702234 427676 702607
rect 427636 702228 427688 702234
rect 427636 702170 427688 702176
rect 437216 701692 437244 703394
rect 447692 703316 447744 703322
rect 447692 703258 447744 703264
rect 447704 701692 447732 703258
rect 458180 703248 458232 703254
rect 458180 703190 458232 703196
rect 458192 701692 458220 703190
rect 419658 701134 419764 701162
rect 419736 701078 419764 701134
rect 422864 701134 423154 701162
rect 429856 701134 430146 701162
rect 433352 701134 433642 701162
rect 440344 701134 440726 701162
rect 443840 701134 444222 701162
rect 450832 701134 451214 701162
rect 454328 701134 454710 701162
rect 461504 701134 461794 701162
rect 422864 701078 422892 701134
rect 429856 701078 429884 701134
rect 433352 701078 433380 701134
rect 440344 701078 440372 701134
rect 443840 701078 443868 701134
rect 450832 701078 450860 701134
rect 454328 701078 454356 701134
rect 461504 701078 461532 701134
rect 462332 701078 462360 703520
rect 468760 703180 468812 703186
rect 468760 703122 468812 703128
rect 468772 701692 468800 703122
rect 475752 702364 475804 702370
rect 475752 702306 475804 702312
rect 472256 702296 472308 702302
rect 472256 702238 472308 702244
rect 472268 701692 472296 702238
rect 475764 701692 475792 702306
rect 465092 701134 465290 701162
rect 465092 701078 465120 701134
rect 478524 701078 478552 703520
rect 479248 703112 479300 703118
rect 479248 703054 479300 703060
rect 479260 701692 479288 703054
rect 489828 703044 489880 703050
rect 489828 702986 489880 702992
rect 486332 702432 486384 702438
rect 486332 702374 486384 702380
rect 486344 701692 486372 702374
rect 489840 701692 489868 702986
rect 494808 702817 494836 703520
rect 500316 702976 500368 702982
rect 500316 702918 500368 702924
rect 494794 702808 494850 702817
rect 494794 702743 494850 702752
rect 496910 701720 496966 701729
rect 496846 701678 496910 701706
rect 500328 701692 500356 702918
rect 514114 701856 514170 701865
rect 514114 701791 514170 701800
rect 514128 701706 514156 701791
rect 514128 701678 514418 701706
rect 496910 701655 496966 701664
rect 492954 701584 493010 701593
rect 503626 701584 503682 701593
rect 493010 701542 493350 701570
rect 492954 701519 493010 701528
rect 503682 701542 503838 701570
rect 503626 701519 503682 701528
rect 506938 701448 506994 701457
rect 517610 701448 517666 701457
rect 506994 701406 507334 701434
rect 506938 701383 506994 701392
rect 517666 701406 517914 701434
rect 517610 701383 517666 701392
rect 524602 701312 524658 701321
rect 482480 701282 482770 701298
rect 482468 701276 482770 701282
rect 482520 701270 482770 701276
rect 524658 701270 524906 701298
rect 524602 701247 524658 701256
rect 482468 701218 482520 701224
rect 527192 701185 527220 703520
rect 543476 703390 543504 703520
rect 543464 703384 543516 703390
rect 543464 703326 543516 703332
rect 542452 702704 542504 702710
rect 542452 702646 542504 702652
rect 538954 702264 539010 702273
rect 538954 702199 539010 702208
rect 538968 701692 538996 702199
rect 542464 701692 542492 702646
rect 552952 701692 552980 703734
rect 559626 703520 559738 704960
rect 563520 703724 563572 703730
rect 563520 703666 563572 703672
rect 559668 702545 559696 703520
rect 559654 702536 559710 702545
rect 559654 702471 559710 702480
rect 556436 702092 556488 702098
rect 556436 702034 556488 702040
rect 556448 701692 556476 702034
rect 563532 701692 563560 703666
rect 575818 703520 575930 704960
rect 577044 703520 577096 703526
rect 577042 703488 577044 703497
rect 577096 703488 577098 703497
rect 577042 703423 577098 703432
rect 582470 702128 582526 702137
rect 582470 702063 582526 702072
rect 532240 701208 532292 701214
rect 510710 701176 510766 701185
rect 521106 701176 521162 701185
rect 510766 701134 510922 701162
rect 510710 701111 510766 701120
rect 527178 701176 527234 701185
rect 521162 701134 521410 701162
rect 521106 701111 521162 701120
rect 527178 701111 527234 701120
rect 528190 701176 528246 701185
rect 531962 701176 532018 701185
rect 528246 701134 528402 701162
rect 531898 701134 531962 701162
rect 528190 701111 528246 701120
rect 531962 701111 532018 701120
rect 532238 701176 532240 701185
rect 535552 701208 535604 701214
rect 532292 701176 532294 701185
rect 535486 701156 535552 701162
rect 535486 701150 535604 701156
rect 545578 701176 545634 701185
rect 535486 701134 535592 701150
rect 532238 701111 532294 701120
rect 549718 701176 549774 701185
rect 545634 701134 545974 701162
rect 549470 701134 549718 701162
rect 545578 701111 545634 701120
rect 549718 701111 549774 701120
rect 559838 701176 559894 701185
rect 570234 701176 570290 701185
rect 559894 701134 560050 701162
rect 566752 701134 567042 701162
rect 559838 701111 559894 701120
rect 566752 701078 566780 701134
rect 573730 701176 573786 701185
rect 570290 701134 570538 701162
rect 570234 701111 570290 701120
rect 581090 701176 581146 701185
rect 573786 701134 574034 701162
rect 577530 701134 577912 701162
rect 581026 701134 581090 701162
rect 573730 701111 573786 701120
rect 577884 701078 577912 701134
rect 581090 701111 581146 701120
rect 184204 701072 184256 701078
rect 184204 701014 184256 701020
rect 202788 701072 202840 701078
rect 202788 701014 202840 701020
rect 262036 701072 262088 701078
rect 262036 701014 262088 701020
rect 265624 701072 265676 701078
rect 265624 701014 265676 701020
rect 267648 701072 267700 701078
rect 267648 701014 267700 701020
rect 283840 701072 283892 701078
rect 283840 701014 283892 701020
rect 318248 701072 318300 701078
rect 318248 701014 318300 701020
rect 332508 701072 332560 701078
rect 332508 701014 332560 701020
rect 333244 701072 333296 701078
rect 333244 701014 333296 701020
rect 349068 701072 349120 701078
rect 349068 701014 349120 701020
rect 356704 701072 356756 701078
rect 356704 701014 356756 701020
rect 360108 701072 360160 701078
rect 360108 701014 360160 701020
rect 398196 701072 398248 701078
rect 398196 701014 398248 701020
rect 401692 701072 401744 701078
rect 401692 701014 401744 701020
rect 404360 701072 404412 701078
rect 404360 701014 404412 701020
rect 419724 701072 419776 701078
rect 419724 701014 419776 701020
rect 422852 701072 422904 701078
rect 422852 701014 422904 701020
rect 429844 701072 429896 701078
rect 429844 701014 429896 701020
rect 433340 701072 433392 701078
rect 433340 701014 433392 701020
rect 440332 701072 440384 701078
rect 440332 701014 440384 701020
rect 443828 701072 443880 701078
rect 443828 701014 443880 701020
rect 450820 701072 450872 701078
rect 450820 701014 450872 701020
rect 454316 701072 454368 701078
rect 454316 701014 454368 701020
rect 461492 701072 461544 701078
rect 461492 701014 461544 701020
rect 462320 701072 462372 701078
rect 462320 701014 462372 701020
rect 465080 701072 465132 701078
rect 465080 701014 465132 701020
rect 478512 701072 478564 701078
rect 478512 701014 478564 701020
rect 566740 701072 566792 701078
rect 566740 701014 566792 701020
rect 577872 701072 577924 701078
rect 577872 701014 577924 701020
rect 580264 302456 580316 302462
rect 580264 302398 580316 302404
rect 183204 299538 183232 301852
rect 183664 301838 183954 301866
rect 184400 301838 184782 301866
rect 184952 301838 185610 301866
rect 183192 299532 183244 299538
rect 183192 299474 183244 299480
rect 183560 299532 183612 299538
rect 183560 299474 183612 299480
rect 183100 46912 183152 46918
rect 183100 46854 183152 46860
rect 183468 10736 183520 10742
rect 183468 10678 183520 10684
rect 182180 4888 182232 4894
rect 182180 4830 182232 4836
rect 183480 3534 183508 10678
rect 183572 4962 183600 299474
rect 183560 4956 183612 4962
rect 183560 4898 183612 4904
rect 183664 4826 183692 301838
rect 184400 299538 184428 301838
rect 184388 299532 184440 299538
rect 184388 299474 184440 299480
rect 184952 6186 184980 301838
rect 186136 10668 186188 10674
rect 186136 10610 186188 10616
rect 184940 6180 184992 6186
rect 184940 6122 184992 6128
rect 183744 5772 183796 5778
rect 183744 5714 183796 5720
rect 183652 4820 183704 4826
rect 183652 4762 183704 4768
rect 181444 3528 181496 3534
rect 181444 3470 181496 3476
rect 182088 3528 182140 3534
rect 182088 3470 182140 3476
rect 182548 3528 182600 3534
rect 182548 3470 182600 3476
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 181456 480 181484 3470
rect 182560 480 182588 3470
rect 183756 480 183784 5714
rect 184940 4820 184992 4826
rect 184940 4762 184992 4768
rect 184952 480 184980 4762
rect 186148 480 186176 10610
rect 186424 3466 186452 301852
rect 187252 298790 187280 301852
rect 187712 301838 188002 301866
rect 188172 301838 188830 301866
rect 189184 301838 189658 301866
rect 187240 298784 187292 298790
rect 187240 298726 187292 298732
rect 187332 6180 187384 6186
rect 187332 6122 187384 6128
rect 186412 3460 186464 3466
rect 186412 3402 186464 3408
rect 187344 480 187372 6122
rect 187712 5030 187740 301838
rect 188172 296714 188200 301838
rect 187804 296686 188200 296714
rect 187804 6254 187832 296686
rect 188988 12096 189040 12102
rect 188988 12038 189040 12044
rect 187792 6248 187844 6254
rect 187792 6190 187844 6196
rect 187700 5024 187752 5030
rect 187700 4966 187752 4972
rect 189000 3534 189028 12038
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 188988 3528 189040 3534
rect 188988 3470 189040 3476
rect 188540 480 188568 3470
rect 189184 2854 189212 301838
rect 190368 10804 190420 10810
rect 190368 10746 190420 10752
rect 190380 3466 190408 10746
rect 190472 3534 190500 301852
rect 190564 301838 191314 301866
rect 190564 5098 190592 301838
rect 192128 297430 192156 301852
rect 192864 298926 192892 301852
rect 192852 298920 192904 298926
rect 192852 298862 192904 298868
rect 193692 298858 193720 301852
rect 193876 301838 194534 301866
rect 194612 301838 195362 301866
rect 196084 301838 196190 301866
rect 196544 301838 196926 301866
rect 197372 301838 197754 301866
rect 197832 301838 198582 301866
rect 193680 298852 193732 298858
rect 193680 298794 193732 298800
rect 192116 297424 192168 297430
rect 192116 297366 192168 297372
rect 193876 296714 193904 301838
rect 193324 296686 193904 296714
rect 190828 6248 190880 6254
rect 190828 6190 190880 6196
rect 190552 5092 190604 5098
rect 190552 5034 190604 5040
rect 190460 3528 190512 3534
rect 190460 3470 190512 3476
rect 189724 3460 189776 3466
rect 189724 3402 189776 3408
rect 190368 3460 190420 3466
rect 190368 3402 190420 3408
rect 189172 2848 189224 2854
rect 189172 2790 189224 2796
rect 189736 480 189764 3402
rect 190840 480 190868 6190
rect 193324 5234 193352 296686
rect 194612 19990 194640 301838
rect 195980 299192 196032 299198
rect 195980 299134 196032 299140
rect 194600 19984 194652 19990
rect 194600 19926 194652 19932
rect 195888 17264 195940 17270
rect 195888 17206 195940 17212
rect 194508 11008 194560 11014
rect 194508 10950 194560 10956
rect 194416 5704 194468 5710
rect 194416 5646 194468 5652
rect 193312 5228 193364 5234
rect 193312 5170 193364 5176
rect 192024 4888 192076 4894
rect 192024 4830 192076 4836
rect 192036 480 192064 4830
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 193232 480 193260 3470
rect 194428 480 194456 5646
rect 194520 3534 194548 10950
rect 195900 6914 195928 17206
rect 195624 6886 195928 6914
rect 194508 3528 194560 3534
rect 194508 3470 194560 3476
rect 195624 480 195652 6886
rect 195992 3738 196020 299134
rect 195980 3732 196032 3738
rect 195980 3674 196032 3680
rect 196084 3670 196112 301838
rect 196544 299198 196572 301838
rect 196532 299192 196584 299198
rect 196532 299134 196584 299140
rect 197268 12232 197320 12238
rect 197268 12174 197320 12180
rect 196072 3664 196124 3670
rect 196072 3606 196124 3612
rect 197280 3534 197308 12174
rect 197372 5166 197400 301838
rect 197832 296714 197860 301838
rect 199396 298926 199424 301852
rect 200224 298994 200252 301852
rect 200316 301838 201066 301866
rect 201604 301838 201802 301866
rect 202248 301838 202630 301866
rect 202892 301838 203458 301866
rect 204286 301838 204392 301866
rect 200212 298988 200264 298994
rect 200212 298930 200264 298936
rect 199384 298920 199436 298926
rect 199384 298862 199436 298868
rect 200316 296714 200344 301838
rect 201500 299192 201552 299198
rect 201500 299134 201552 299140
rect 197464 296686 197860 296714
rect 200224 296686 200344 296714
rect 197464 296002 197492 296686
rect 197452 295996 197504 296002
rect 197452 295938 197504 295944
rect 200028 13116 200080 13122
rect 200028 13058 200080 13064
rect 197912 5636 197964 5642
rect 197912 5578 197964 5584
rect 197360 5160 197412 5166
rect 197360 5102 197412 5108
rect 196808 3528 196860 3534
rect 196808 3470 196860 3476
rect 197268 3528 197320 3534
rect 197268 3470 197320 3476
rect 196820 480 196848 3470
rect 197924 480 197952 5578
rect 200040 3466 200068 13058
rect 200224 5302 200252 296686
rect 201512 16574 201540 299134
rect 201604 294642 201632 301838
rect 202248 299198 202276 301838
rect 202236 299192 202288 299198
rect 202236 299134 202288 299140
rect 201592 294636 201644 294642
rect 201592 294578 201644 294584
rect 201512 16546 201632 16574
rect 200212 5296 200264 5302
rect 200212 5238 200264 5244
rect 201500 5092 201552 5098
rect 201500 5034 201552 5040
rect 199108 3460 199160 3466
rect 199108 3402 199160 3408
rect 200028 3460 200080 3466
rect 200028 3402 200080 3408
rect 200304 3460 200356 3466
rect 200304 3402 200356 3408
rect 199120 480 199148 3402
rect 200316 480 200344 3402
rect 201512 480 201540 5034
rect 201604 3738 201632 16546
rect 202892 5370 202920 301838
rect 204364 39370 204392 301838
rect 205100 299062 205128 301852
rect 205652 301838 205850 301866
rect 206296 301838 206678 301866
rect 207032 301838 207506 301866
rect 207584 301838 208334 301866
rect 208412 301838 209162 301866
rect 205088 299056 205140 299062
rect 205088 298998 205140 299004
rect 204352 39364 204404 39370
rect 204352 39306 204404 39312
rect 205652 5438 205680 301838
rect 206296 296714 206324 301838
rect 205744 296686 206324 296714
rect 205744 294710 205772 296686
rect 205732 294704 205784 294710
rect 205732 294646 205784 294652
rect 206192 8832 206244 8838
rect 206192 8774 206244 8780
rect 205640 5432 205692 5438
rect 205640 5374 205692 5380
rect 202880 5364 202932 5370
rect 202880 5306 202932 5312
rect 205088 5024 205140 5030
rect 205088 4966 205140 4972
rect 202696 4956 202748 4962
rect 202696 4898 202748 4904
rect 201592 3732 201644 3738
rect 201592 3674 201644 3680
rect 202708 480 202736 4898
rect 203892 3596 203944 3602
rect 203892 3538 203944 3544
rect 203904 480 203932 3538
rect 205100 480 205128 4966
rect 206204 480 206232 8774
rect 207032 3874 207060 301838
rect 207584 296714 207612 301838
rect 207124 296686 207612 296714
rect 207124 7614 207152 296686
rect 208412 296070 208440 301838
rect 209976 299130 210004 301852
rect 210160 301838 210726 301866
rect 209964 299124 210016 299130
rect 209964 299066 210016 299072
rect 210160 296714 210188 301838
rect 210424 298852 210476 298858
rect 210424 298794 210476 298800
rect 209884 296686 210188 296714
rect 208400 296064 208452 296070
rect 208400 296006 208452 296012
rect 209688 295996 209740 296002
rect 209688 295938 209740 295944
rect 207112 7608 207164 7614
rect 207112 7550 207164 7556
rect 207020 3868 207072 3874
rect 207020 3810 207072 3816
rect 207388 3664 207440 3670
rect 207388 3606 207440 3612
rect 207400 480 207428 3606
rect 209700 3534 209728 295938
rect 209780 8696 209832 8702
rect 209780 8638 209832 8644
rect 208584 3528 208636 3534
rect 208584 3470 208636 3476
rect 209688 3528 209740 3534
rect 209688 3470 209740 3476
rect 208596 480 208624 3470
rect 209792 480 209820 8638
rect 209884 7682 209912 296686
rect 209872 7676 209924 7682
rect 209872 7618 209924 7624
rect 210436 4010 210464 298794
rect 211540 297498 211568 301852
rect 211724 301838 212382 301866
rect 212552 301838 213210 301866
rect 211528 297492 211580 297498
rect 211528 297434 211580 297440
rect 211724 296714 211752 301838
rect 211804 298920 211856 298926
rect 211804 298862 211856 298868
rect 211172 296686 211752 296714
rect 210424 4004 210476 4010
rect 210424 3946 210476 3952
rect 211172 3806 211200 296686
rect 211816 3942 211844 298862
rect 212552 7750 212580 301838
rect 214024 296138 214052 301852
rect 214760 299266 214788 301852
rect 215312 301838 215602 301866
rect 215680 301838 216430 301866
rect 214748 299260 214800 299266
rect 214748 299202 214800 299208
rect 214564 298988 214616 298994
rect 214564 298930 214616 298936
rect 214012 296132 214064 296138
rect 214012 296074 214064 296080
rect 213368 8764 213420 8770
rect 213368 8706 213420 8712
rect 212540 7744 212592 7750
rect 212540 7686 212592 7692
rect 212540 5160 212592 5166
rect 212540 5102 212592 5108
rect 211804 3936 211856 3942
rect 211804 3878 211856 3884
rect 211160 3800 211212 3806
rect 211160 3742 211212 3748
rect 210976 3732 211028 3738
rect 210976 3674 211028 3680
rect 210988 480 211016 3674
rect 212552 2802 212580 5102
rect 212184 2774 212580 2802
rect 212184 480 212212 2774
rect 213380 480 213408 8706
rect 214472 3800 214524 3806
rect 214472 3742 214524 3748
rect 214484 480 214512 3742
rect 214576 3398 214604 298930
rect 214656 298784 214708 298790
rect 214656 298726 214708 298732
rect 214668 4146 214696 298726
rect 215312 5506 215340 301838
rect 215680 296714 215708 301838
rect 217244 298382 217272 301852
rect 217324 299124 217376 299130
rect 217324 299066 217376 299072
rect 217232 298376 217284 298382
rect 217232 298318 217284 298324
rect 215404 296686 215708 296714
rect 215404 7818 215432 296686
rect 216864 8628 216916 8634
rect 216864 8570 216916 8576
rect 215392 7812 215444 7818
rect 215392 7754 215444 7760
rect 215300 5500 215352 5506
rect 215300 5442 215352 5448
rect 215668 5228 215720 5234
rect 215668 5170 215720 5176
rect 214656 4140 214708 4146
rect 214656 4082 214708 4088
rect 214564 3392 214616 3398
rect 214564 3334 214616 3340
rect 215680 480 215708 5170
rect 216876 480 216904 8570
rect 217336 3330 217364 299066
rect 218072 4758 218100 301852
rect 218164 301838 218914 301866
rect 218164 7886 218192 301838
rect 219636 298858 219664 301852
rect 219728 301838 220478 301866
rect 220924 301838 221306 301866
rect 219624 298852 219676 298858
rect 219624 298794 219676 298800
rect 219728 296714 219756 301838
rect 220084 299192 220136 299198
rect 220084 299134 220136 299140
rect 219544 296686 219756 296714
rect 218152 7880 218204 7886
rect 218152 7822 218204 7828
rect 218060 4752 218112 4758
rect 218060 4694 218112 4700
rect 219544 4690 219572 296686
rect 219532 4684 219584 4690
rect 219532 4626 219584 4632
rect 219256 4004 219308 4010
rect 219256 3946 219308 3952
rect 218060 3528 218112 3534
rect 218060 3470 218112 3476
rect 217324 3324 217376 3330
rect 217324 3266 217376 3272
rect 218072 480 218100 3470
rect 219268 480 219296 3946
rect 220096 3262 220124 299134
rect 220452 8560 220504 8566
rect 220452 8502 220504 8508
rect 220084 3256 220136 3262
rect 220084 3198 220136 3204
rect 220464 480 220492 8502
rect 220924 7954 220952 301838
rect 222120 298450 222148 301852
rect 222212 301838 222962 301866
rect 222108 298444 222160 298450
rect 222108 298386 222160 298392
rect 221464 298376 221516 298382
rect 221464 298318 221516 298324
rect 220912 7948 220964 7954
rect 220912 7890 220964 7896
rect 221476 3194 221504 298318
rect 222212 4554 222240 301838
rect 223488 296064 223540 296070
rect 223488 296006 223540 296012
rect 222200 4548 222252 4554
rect 222200 4490 222252 4496
rect 221556 4072 221608 4078
rect 221556 4014 221608 4020
rect 221464 3188 221516 3194
rect 221464 3130 221516 3136
rect 221568 480 221596 4014
rect 223500 3398 223528 296006
rect 223684 8022 223712 301852
rect 224512 298926 224540 301852
rect 224972 301838 225354 301866
rect 225432 301838 226182 301866
rect 224500 298920 224552 298926
rect 224500 298862 224552 298868
rect 224224 298852 224276 298858
rect 224224 298794 224276 298800
rect 223948 8424 224000 8430
rect 223948 8366 224000 8372
rect 223672 8016 223724 8022
rect 223672 7958 223724 7964
rect 222752 3392 222804 3398
rect 222752 3334 222804 3340
rect 223488 3392 223540 3398
rect 223488 3334 223540 3340
rect 222764 480 222792 3334
rect 223960 480 223988 8366
rect 224236 3126 224264 298794
rect 224972 4622 225000 301838
rect 225432 296714 225460 301838
rect 226996 298518 227024 301852
rect 227732 301838 227838 301866
rect 228008 301838 228574 301866
rect 227076 299056 227128 299062
rect 227076 298998 227128 299004
rect 226984 298512 227036 298518
rect 226984 298454 227036 298460
rect 227088 296714 227116 298998
rect 225064 296686 225460 296714
rect 226996 296686 227116 296714
rect 225064 8090 225092 296686
rect 225052 8084 225104 8090
rect 225052 8026 225104 8032
rect 224960 4616 225012 4622
rect 224960 4558 225012 4564
rect 226340 4140 226392 4146
rect 226340 4082 226392 4088
rect 225144 3936 225196 3942
rect 225144 3878 225196 3884
rect 224224 3120 224276 3126
rect 224224 3062 224276 3068
rect 225156 480 225184 3878
rect 226352 480 226380 4082
rect 226996 3058 227024 296686
rect 227536 8492 227588 8498
rect 227536 8434 227588 8440
rect 226984 3052 227036 3058
rect 226984 2994 227036 3000
rect 227548 480 227576 8434
rect 227732 4486 227760 301838
rect 228008 296714 228036 301838
rect 229388 298790 229416 301852
rect 229480 301838 230230 301866
rect 230492 301838 231058 301866
rect 229376 298784 229428 298790
rect 229376 298726 229428 298732
rect 229480 296714 229508 301838
rect 227824 296686 228036 296714
rect 229204 296686 229508 296714
rect 227824 8158 227852 296686
rect 227812 8152 227864 8158
rect 227812 8094 227864 8100
rect 227720 4480 227772 4486
rect 227720 4422 227772 4428
rect 229204 4350 229232 296686
rect 230492 8226 230520 301838
rect 230572 298784 230624 298790
rect 230572 298726 230624 298732
rect 230584 294914 230612 298726
rect 231872 298314 231900 301852
rect 231964 301838 232622 301866
rect 233344 301838 233450 301866
rect 231860 298308 231912 298314
rect 231860 298250 231912 298256
rect 230572 294908 230624 294914
rect 230572 294850 230624 294856
rect 231768 294636 231820 294642
rect 231768 294578 231820 294584
rect 230480 8220 230532 8226
rect 230480 8162 230532 8168
rect 231400 5296 231452 5302
rect 231400 5238 231452 5244
rect 229192 4344 229244 4350
rect 229192 4286 229244 4292
rect 231032 3460 231084 3466
rect 231032 3402 231084 3408
rect 228732 3324 228784 3330
rect 228732 3266 228784 3272
rect 228744 480 228772 3266
rect 229836 2848 229888 2854
rect 229836 2790 229888 2796
rect 229848 480 229876 2790
rect 231044 480 231072 3402
rect 231412 2854 231440 5238
rect 231780 3466 231808 294578
rect 231964 4418 231992 301838
rect 232504 299260 232556 299266
rect 232504 299202 232556 299208
rect 231952 4412 232004 4418
rect 231952 4354 232004 4360
rect 231768 3460 231820 3466
rect 231768 3402 231820 3408
rect 232228 3460 232280 3466
rect 232228 3402 232280 3408
rect 231400 2848 231452 2854
rect 231400 2790 231452 2796
rect 232240 480 232268 3402
rect 232516 2990 232544 299202
rect 233344 8294 233372 301838
rect 234264 298994 234292 301852
rect 234632 301838 235106 301866
rect 235184 301838 235934 301866
rect 234252 298988 234304 298994
rect 234252 298930 234304 298936
rect 234528 298988 234580 298994
rect 234528 298930 234580 298936
rect 234540 298178 234568 298930
rect 233884 298172 233936 298178
rect 233884 298114 233936 298120
rect 234528 298172 234580 298178
rect 234528 298114 234580 298120
rect 233332 8288 233384 8294
rect 233332 8230 233384 8236
rect 233424 7676 233476 7682
rect 233424 7618 233476 7624
rect 232504 2984 232556 2990
rect 232504 2926 232556 2932
rect 233436 480 233464 7618
rect 233896 2922 233924 298114
rect 234632 4282 234660 301838
rect 235184 296714 235212 301838
rect 236748 298246 236776 301852
rect 237392 301838 237498 301866
rect 237944 301838 238326 301866
rect 236736 298240 236788 298246
rect 236736 298182 236788 298188
rect 234724 296686 235212 296714
rect 234724 7546 234752 296686
rect 237012 7608 237064 7614
rect 237012 7550 237064 7556
rect 234712 7540 234764 7546
rect 234712 7482 234764 7488
rect 234620 4276 234672 4282
rect 234620 4218 234672 4224
rect 234620 3868 234672 3874
rect 234620 3810 234672 3816
rect 233884 2916 233936 2922
rect 233884 2858 233936 2864
rect 234632 480 234660 3810
rect 235816 3256 235868 3262
rect 235816 3198 235868 3204
rect 235828 480 235856 3198
rect 237024 480 237052 7550
rect 237392 6322 237420 301838
rect 237944 296714 237972 301838
rect 239140 299130 239168 301852
rect 239232 301838 239982 301866
rect 239128 299124 239180 299130
rect 239128 299066 239180 299072
rect 239232 296714 239260 301838
rect 240796 297566 240824 301852
rect 240874 300248 240930 300257
rect 240874 300183 240930 300192
rect 240784 297560 240836 297566
rect 240784 297502 240836 297508
rect 237484 296686 237972 296714
rect 238864 296686 239260 296714
rect 237484 14482 237512 296686
rect 237472 14476 237524 14482
rect 237472 14418 237524 14424
rect 238024 14476 238076 14482
rect 238024 14418 238076 14424
rect 237380 6316 237432 6322
rect 237380 6258 237432 6264
rect 238036 3330 238064 14418
rect 238864 6390 238892 296686
rect 240784 296132 240836 296138
rect 240784 296074 240836 296080
rect 240508 7744 240560 7750
rect 240508 7686 240560 7692
rect 238852 6384 238904 6390
rect 238852 6326 238904 6332
rect 238116 3392 238168 3398
rect 238116 3334 238168 3340
rect 238024 3324 238076 3330
rect 238024 3266 238076 3272
rect 238128 480 238156 3334
rect 239312 3188 239364 3194
rect 239312 3130 239364 3136
rect 239324 480 239352 3130
rect 240520 480 240548 7686
rect 240796 3874 240824 296074
rect 240888 139398 240916 300183
rect 241624 299198 241652 301852
rect 241900 301838 242374 301866
rect 241612 299192 241664 299198
rect 241612 299134 241664 299140
rect 241900 296714 241928 301838
rect 243188 297634 243216 301852
rect 244016 299334 244044 301852
rect 244292 301838 244858 301866
rect 244004 299328 244056 299334
rect 244004 299270 244056 299276
rect 243176 297628 243228 297634
rect 243176 297570 243228 297576
rect 242164 297424 242216 297430
rect 242164 297366 242216 297372
rect 241624 296686 241928 296714
rect 240968 140072 241020 140078
rect 240968 140014 241020 140020
rect 240876 139392 240928 139398
rect 240876 139334 240928 139340
rect 240784 3868 240836 3874
rect 240784 3810 240836 3816
rect 240980 3262 241008 140014
rect 241624 6458 241652 296686
rect 241612 6452 241664 6458
rect 241612 6394 241664 6400
rect 241704 3460 241756 3466
rect 241704 3402 241756 3408
rect 240968 3256 241020 3262
rect 240968 3198 241020 3204
rect 241716 480 241744 3402
rect 242176 3330 242204 297366
rect 244096 7812 244148 7818
rect 244096 7754 244148 7760
rect 242164 3324 242216 3330
rect 242164 3266 242216 3272
rect 242900 3256 242952 3262
rect 242900 3198 242952 3204
rect 242912 480 242940 3198
rect 244108 480 244136 7754
rect 244292 6526 244320 301838
rect 245672 297702 245700 301852
rect 246408 298858 246436 301852
rect 247144 301838 247250 301866
rect 246948 299328 247000 299334
rect 246948 299270 247000 299276
rect 246488 299192 246540 299198
rect 246488 299134 246540 299140
rect 246396 298852 246448 298858
rect 246396 298794 246448 298800
rect 245660 297696 245712 297702
rect 245660 297638 245712 297644
rect 244924 297492 244976 297498
rect 244924 297434 244976 297440
rect 244280 6520 244332 6526
rect 244280 6462 244332 6468
rect 244936 3194 244964 297434
rect 246304 297152 246356 297158
rect 246304 297094 246356 297100
rect 246316 3534 246344 297094
rect 246500 296714 246528 299134
rect 246408 296686 246528 296714
rect 246408 10266 246436 296686
rect 246960 296206 246988 299270
rect 246948 296200 247000 296206
rect 246948 296142 247000 296148
rect 246396 10260 246448 10266
rect 246396 10202 246448 10208
rect 247144 6594 247172 301838
rect 248064 299334 248092 301852
rect 248052 299328 248104 299334
rect 248052 299270 248104 299276
rect 248892 298722 248920 301852
rect 248984 301838 249734 301866
rect 249812 301838 250562 301866
rect 248880 298716 248932 298722
rect 248880 298658 248932 298664
rect 248984 296714 249012 301838
rect 249064 298852 249116 298858
rect 249064 298794 249116 298800
rect 248524 296686 249012 296714
rect 247592 7880 247644 7886
rect 247592 7822 247644 7828
rect 247132 6588 247184 6594
rect 247132 6530 247184 6536
rect 246304 3528 246356 3534
rect 246304 3470 246356 3476
rect 246396 3324 246448 3330
rect 246396 3266 246448 3272
rect 244924 3188 244976 3194
rect 244924 3130 244976 3136
rect 245200 3188 245252 3194
rect 245200 3130 245252 3136
rect 245212 480 245240 3130
rect 246408 480 246436 3266
rect 247604 480 247632 7822
rect 248524 6662 248552 296686
rect 248512 6656 248564 6662
rect 248512 6598 248564 6604
rect 248788 3596 248840 3602
rect 248788 3538 248840 3544
rect 248800 480 248828 3538
rect 249076 3398 249104 298794
rect 249812 296274 249840 301838
rect 251284 298926 251312 301852
rect 251376 301838 252126 301866
rect 251272 298920 251324 298926
rect 251272 298862 251324 298868
rect 250536 298512 250588 298518
rect 250536 298454 250588 298460
rect 250444 297084 250496 297090
rect 250444 297026 250496 297032
rect 249800 296268 249852 296274
rect 249800 296210 249852 296216
rect 250456 6914 250484 297026
rect 250548 13190 250576 298454
rect 251376 296714 251404 301838
rect 251732 298716 251784 298722
rect 251732 298658 251784 298664
rect 251284 296686 251404 296714
rect 250536 13184 250588 13190
rect 250536 13126 250588 13132
rect 251088 12164 251140 12170
rect 251088 12106 251140 12112
rect 249904 6886 250484 6914
rect 249904 3534 249932 6886
rect 251100 3534 251128 12106
rect 251180 7948 251232 7954
rect 251180 7890 251232 7896
rect 249892 3528 249944 3534
rect 249892 3470 249944 3476
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 251088 3528 251140 3534
rect 251088 3470 251140 3476
rect 249064 3392 249116 3398
rect 249064 3334 249116 3340
rect 249996 480 250024 3470
rect 251192 480 251220 7890
rect 251284 7478 251312 296686
rect 251744 294846 251772 298658
rect 252940 297770 252968 301852
rect 253768 299402 253796 301852
rect 253952 301838 254610 301866
rect 255346 301838 255452 301866
rect 253756 299396 253808 299402
rect 253756 299338 253808 299344
rect 253296 299328 253348 299334
rect 253296 299270 253348 299276
rect 253204 299124 253256 299130
rect 253204 299066 253256 299072
rect 252928 297764 252980 297770
rect 252928 297706 252980 297712
rect 251824 295792 251876 295798
rect 251824 295734 251876 295740
rect 251732 294840 251784 294846
rect 251732 294782 251784 294788
rect 251272 7472 251324 7478
rect 251272 7414 251324 7420
rect 251836 4010 251864 295734
rect 253216 10878 253244 299066
rect 253308 12034 253336 299270
rect 253388 13184 253440 13190
rect 253388 13126 253440 13132
rect 253296 12028 253348 12034
rect 253296 11970 253348 11976
rect 253204 10872 253256 10878
rect 253204 10814 253256 10820
rect 253400 4078 253428 13126
rect 253848 10872 253900 10878
rect 253848 10814 253900 10820
rect 253388 4072 253440 4078
rect 253388 4014 253440 4020
rect 251824 4004 251876 4010
rect 251824 3946 251876 3952
rect 252376 3392 252428 3398
rect 252376 3334 252428 3340
rect 252388 480 252416 3334
rect 253492 598 253704 626
rect 253492 480 253520 598
rect 253676 490 253704 598
rect 253860 490 253888 10814
rect 253952 8974 253980 301838
rect 255424 296342 255452 301838
rect 256160 299470 256188 301852
rect 256712 301838 257002 301866
rect 256148 299464 256200 299470
rect 256148 299406 256200 299412
rect 255964 298920 256016 298926
rect 255964 298862 256016 298868
rect 255412 296336 255464 296342
rect 255412 296278 255464 296284
rect 253940 8968 253992 8974
rect 253940 8910 253992 8916
rect 254676 4004 254728 4010
rect 254676 3946 254728 3952
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 253676 462 253888 490
rect 254688 480 254716 3946
rect 255872 3596 255924 3602
rect 255872 3538 255924 3544
rect 255884 480 255912 3538
rect 255976 3194 256004 298862
rect 256056 295860 256108 295866
rect 256056 295802 256108 295808
rect 256068 4146 256096 295802
rect 256712 9110 256740 301838
rect 257816 297838 257844 301852
rect 258080 299464 258132 299470
rect 258080 299406 258132 299412
rect 257804 297832 257856 297838
rect 257804 297774 257856 297780
rect 258092 294778 258120 299406
rect 258644 299062 258672 301852
rect 258632 299056 258684 299062
rect 258632 298998 258684 299004
rect 258816 298512 258868 298518
rect 258816 298454 258868 298460
rect 258724 297016 258776 297022
rect 258724 296958 258776 296964
rect 258080 294772 258132 294778
rect 258080 294714 258132 294720
rect 256700 9104 256752 9110
rect 256700 9046 256752 9052
rect 258736 4146 258764 296958
rect 258828 10946 258856 298454
rect 258816 10940 258868 10946
rect 258816 10882 258868 10888
rect 259368 10940 259420 10946
rect 259368 10882 259420 10888
rect 256056 4140 256108 4146
rect 256056 4082 256108 4088
rect 258172 4140 258224 4146
rect 258172 4082 258224 4088
rect 258724 4140 258776 4146
rect 258724 4082 258776 4088
rect 257068 4072 257120 4078
rect 257068 4014 257120 4020
rect 255964 3188 256016 3194
rect 255964 3130 256016 3136
rect 257080 480 257108 4014
rect 258184 3670 258212 4082
rect 259380 3670 259408 10882
rect 259472 9042 259500 301852
rect 259564 301838 260222 301866
rect 259564 296410 259592 301838
rect 261036 298654 261064 301852
rect 261312 301838 261878 301866
rect 261024 298648 261076 298654
rect 261024 298590 261076 298596
rect 260104 297832 260156 297838
rect 260104 297774 260156 297780
rect 259552 296404 259604 296410
rect 259552 296346 259604 296352
rect 259460 9036 259512 9042
rect 259460 8978 259512 8984
rect 259460 4140 259512 4146
rect 259460 4082 259512 4088
rect 258172 3664 258224 3670
rect 258172 3606 258224 3612
rect 258264 3664 258316 3670
rect 258264 3606 258316 3612
rect 259368 3664 259420 3670
rect 259368 3606 259420 3612
rect 258276 480 258304 3606
rect 259472 480 259500 4082
rect 260116 3262 260144 297774
rect 261312 296714 261340 301838
rect 262692 298722 262720 301852
rect 263520 299266 263548 301852
rect 263612 301838 264270 301866
rect 263508 299260 263560 299266
rect 263508 299202 263560 299208
rect 262864 299056 262916 299062
rect 262864 298998 262916 299004
rect 262680 298716 262732 298722
rect 262680 298658 262732 298664
rect 262876 297226 262904 298998
rect 263048 298172 263100 298178
rect 263048 298114 263100 298120
rect 262864 297220 262916 297226
rect 262864 297162 262916 297168
rect 262864 296948 262916 296954
rect 262864 296890 262916 296896
rect 260944 296686 261340 296714
rect 260944 9178 260972 296686
rect 260932 9172 260984 9178
rect 260932 9114 260984 9120
rect 262876 3806 262904 296890
rect 262956 296200 263008 296206
rect 262956 296142 263008 296148
rect 262864 3800 262916 3806
rect 262864 3742 262916 3748
rect 262968 3670 262996 296142
rect 263060 10606 263088 298114
rect 263048 10600 263100 10606
rect 263048 10542 263100 10548
rect 263612 10402 263640 301838
rect 265084 299470 265112 301852
rect 265072 299464 265124 299470
rect 265072 299406 265124 299412
rect 263692 299260 263744 299266
rect 263692 299202 263744 299208
rect 263704 298042 263732 299202
rect 265912 298586 265940 301852
rect 266464 301838 266754 301866
rect 266360 298716 266412 298722
rect 266360 298658 266412 298664
rect 265900 298580 265952 298586
rect 265900 298522 265952 298528
rect 266372 298110 266400 298658
rect 266360 298104 266412 298110
rect 266360 298046 266412 298052
rect 263692 298036 263744 298042
rect 263692 297978 263744 297984
rect 264244 297220 264296 297226
rect 264244 297162 264296 297168
rect 263600 10396 263652 10402
rect 263600 10338 263652 10344
rect 264256 3942 264284 297162
rect 266464 10470 266492 301838
rect 267568 298790 267596 301852
rect 268396 298994 268424 301852
rect 268384 298988 268436 298994
rect 268384 298930 268436 298936
rect 268844 298988 268896 298994
rect 268844 298930 268896 298936
rect 267556 298784 267608 298790
rect 267556 298726 267608 298732
rect 268384 298784 268436 298790
rect 268384 298726 268436 298732
rect 267004 298036 267056 298042
rect 267004 297978 267056 297984
rect 266452 10464 266504 10470
rect 266452 10406 266504 10412
rect 264888 10396 264940 10402
rect 264888 10338 264940 10344
rect 264244 3936 264296 3942
rect 264244 3878 264296 3884
rect 263048 3732 263100 3738
rect 263048 3674 263100 3680
rect 261760 3664 261812 3670
rect 261760 3606 261812 3612
rect 262956 3664 263008 3670
rect 262956 3606 263008 3612
rect 260104 3256 260156 3262
rect 260104 3198 260156 3204
rect 260656 3256 260708 3262
rect 260656 3198 260708 3204
rect 260668 480 260696 3198
rect 261772 480 261800 3606
rect 263060 1850 263088 3674
rect 264900 3670 264928 10338
rect 266544 3936 266596 3942
rect 266544 3878 266596 3884
rect 264152 3664 264204 3670
rect 264152 3606 264204 3612
rect 264888 3664 264940 3670
rect 264888 3606 264940 3612
rect 265348 3664 265400 3670
rect 265348 3606 265400 3612
rect 262968 1822 263088 1850
rect 262968 480 262996 1822
rect 264164 480 264192 3606
rect 265360 480 265388 3606
rect 266556 480 266584 3878
rect 267016 3194 267044 297978
rect 267096 14544 267148 14550
rect 267096 14486 267148 14492
rect 267108 3670 267136 14486
rect 268396 3942 268424 298726
rect 268476 297696 268528 297702
rect 268476 297638 268528 297644
rect 268384 3936 268436 3942
rect 268384 3878 268436 3884
rect 267740 3732 267792 3738
rect 267740 3674 267792 3680
rect 267096 3664 267148 3670
rect 267096 3606 267148 3612
rect 267004 3188 267056 3194
rect 267004 3130 267056 3136
rect 267752 480 267780 3674
rect 268488 3262 268516 297638
rect 268856 297294 268884 298930
rect 269132 298178 269160 301852
rect 269224 301838 269974 301866
rect 270512 301838 270802 301866
rect 269120 298172 269172 298178
rect 269120 298114 269172 298120
rect 268844 297288 268896 297294
rect 268844 297230 268896 297236
rect 269224 6730 269252 301838
rect 269764 297628 269816 297634
rect 269764 297570 269816 297576
rect 269212 6724 269264 6730
rect 269212 6666 269264 6672
rect 269776 3738 269804 297570
rect 269856 10600 269908 10606
rect 269856 10542 269908 10548
rect 269764 3732 269816 3738
rect 269764 3674 269816 3680
rect 269868 3330 269896 10542
rect 270512 7410 270540 301838
rect 271616 297906 271644 301852
rect 271984 301838 272458 301866
rect 271604 297900 271656 297906
rect 271604 297842 271656 297848
rect 271788 297560 271840 297566
rect 271788 297502 271840 297508
rect 271144 14612 271196 14618
rect 271144 14554 271196 14560
rect 270500 7404 270552 7410
rect 270500 7346 270552 7352
rect 271156 4078 271184 14554
rect 271144 4072 271196 4078
rect 271144 4014 271196 4020
rect 270040 3800 270092 3806
rect 270040 3742 270092 3748
rect 269856 3324 269908 3330
rect 269856 3266 269908 3272
rect 268476 3256 268528 3262
rect 268476 3198 268528 3204
rect 268844 3120 268896 3126
rect 268844 3062 268896 3068
rect 268856 480 268884 3062
rect 270052 480 270080 3742
rect 271800 3738 271828 297502
rect 271984 6798 272012 301838
rect 273180 299402 273208 301852
rect 273168 299396 273220 299402
rect 273168 299338 273220 299344
rect 274008 297974 274036 301852
rect 274088 299396 274140 299402
rect 274088 299338 274140 299344
rect 273996 297968 274048 297974
rect 273996 297910 274048 297916
rect 274100 296714 274128 299338
rect 274836 299266 274864 301852
rect 275112 301838 275678 301866
rect 276032 301838 276506 301866
rect 276676 301838 277334 301866
rect 277412 301838 278070 301866
rect 274824 299260 274876 299266
rect 274824 299202 274876 299208
rect 274548 298648 274600 298654
rect 274548 298590 274600 298596
rect 274008 296686 274128 296714
rect 273904 296404 273956 296410
rect 273904 296346 273956 296352
rect 271972 6792 272024 6798
rect 271972 6734 272024 6740
rect 273916 4010 273944 296346
rect 274008 12238 274036 296686
rect 274560 295934 274588 298590
rect 275112 296714 275140 301838
rect 274744 296686 275140 296714
rect 274548 295928 274600 295934
rect 274548 295870 274600 295876
rect 274088 141432 274140 141438
rect 274088 141374 274140 141380
rect 273996 12232 274048 12238
rect 273996 12174 274048 12180
rect 273904 4004 273956 4010
rect 273904 3946 273956 3952
rect 272432 3936 272484 3942
rect 272432 3878 272484 3884
rect 271236 3732 271288 3738
rect 271236 3674 271288 3680
rect 271788 3732 271840 3738
rect 271788 3674 271840 3680
rect 271248 480 271276 3674
rect 272444 480 272472 3878
rect 274100 3874 274128 141374
rect 274744 9246 274772 296686
rect 276032 10538 276060 301838
rect 276676 296714 276704 301838
rect 276124 296686 276704 296714
rect 276124 202162 276152 296686
rect 276112 202156 276164 202162
rect 276112 202098 276164 202104
rect 276664 202156 276716 202162
rect 276664 202098 276716 202104
rect 276020 10532 276072 10538
rect 276020 10474 276072 10480
rect 274732 9240 274784 9246
rect 274732 9182 274784 9188
rect 276020 4004 276072 4010
rect 276020 3946 276072 3952
rect 274088 3868 274140 3874
rect 274088 3810 274140 3816
rect 274824 3324 274876 3330
rect 274824 3266 274876 3272
rect 273628 3256 273680 3262
rect 273628 3198 273680 3204
rect 273640 480 273668 3198
rect 274836 480 274864 3266
rect 276032 480 276060 3946
rect 276676 3126 276704 202098
rect 276756 10464 276808 10470
rect 276756 10406 276808 10412
rect 276768 3330 276796 10406
rect 277412 9314 277440 301838
rect 278884 298722 278912 301852
rect 279712 299062 279740 301852
rect 280264 301838 280554 301866
rect 281000 301838 281382 301866
rect 281552 301838 282118 301866
rect 282946 301838 283052 301866
rect 279700 299056 279752 299062
rect 279700 298998 279752 299004
rect 278872 298716 278924 298722
rect 278872 298658 278924 298664
rect 278044 298580 278096 298586
rect 278044 298522 278096 298528
rect 277400 9308 277452 9314
rect 277400 9250 277452 9256
rect 277124 3800 277176 3806
rect 277124 3742 277176 3748
rect 276756 3324 276808 3330
rect 276756 3266 276808 3272
rect 276664 3120 276716 3126
rect 276664 3062 276716 3068
rect 277136 480 277164 3742
rect 278056 3398 278084 298522
rect 280264 9382 280292 301838
rect 281000 298994 281028 301838
rect 281356 299260 281408 299266
rect 281356 299202 281408 299208
rect 280988 298988 281040 298994
rect 280988 298930 281040 298936
rect 280804 297764 280856 297770
rect 280804 297706 280856 297712
rect 280252 9376 280304 9382
rect 280252 9318 280304 9324
rect 279516 3936 279568 3942
rect 279516 3878 279568 3884
rect 278044 3392 278096 3398
rect 278044 3334 278096 3340
rect 278320 3392 278372 3398
rect 278320 3334 278372 3340
rect 278332 480 278360 3334
rect 279528 480 279556 3878
rect 280816 3398 280844 297706
rect 281368 296546 281396 299202
rect 281356 296540 281408 296546
rect 281356 296482 281408 296488
rect 281552 11762 281580 301838
rect 282184 299056 282236 299062
rect 282184 298998 282236 299004
rect 281540 11756 281592 11762
rect 281540 11698 281592 11704
rect 281908 6316 281960 6322
rect 281908 6258 281960 6264
rect 280804 3392 280856 3398
rect 280804 3334 280856 3340
rect 280712 3120 280764 3126
rect 280712 3062 280764 3068
rect 280724 480 280752 3062
rect 281920 480 281948 6258
rect 282196 3262 282224 298998
rect 283024 9450 283052 301838
rect 283760 299266 283788 301852
rect 283748 299260 283800 299266
rect 283748 299202 283800 299208
rect 284588 298654 284616 301852
rect 284680 301838 285430 301866
rect 285784 301838 286258 301866
rect 286704 301838 286994 301866
rect 287072 301838 287822 301866
rect 288452 301838 288650 301866
rect 288728 301838 289478 301866
rect 289924 301838 290306 301866
rect 284576 298648 284628 298654
rect 284576 298590 284628 298596
rect 284680 296714 284708 301838
rect 285680 299260 285732 299266
rect 285680 299202 285732 299208
rect 284944 298988 284996 298994
rect 284944 298930 284996 298936
rect 284404 296686 284708 296714
rect 284404 9586 284432 296686
rect 284392 9580 284444 9586
rect 284392 9522 284444 9528
rect 283012 9444 283064 9450
rect 283012 9386 283064 9392
rect 284300 3868 284352 3874
rect 284300 3810 284352 3816
rect 283104 3392 283156 3398
rect 283104 3334 283156 3340
rect 282184 3256 282236 3262
rect 282184 3198 282236 3204
rect 283116 480 283144 3334
rect 284312 480 284340 3810
rect 284956 3126 284984 298930
rect 285692 188358 285720 299202
rect 285784 296478 285812 301838
rect 286704 299266 286732 301838
rect 286692 299260 286744 299266
rect 286692 299202 286744 299208
rect 285772 296472 285824 296478
rect 285772 296414 285824 296420
rect 286324 296268 286376 296274
rect 286324 296210 286376 296216
rect 285680 188352 285732 188358
rect 285680 188294 285732 188300
rect 285404 6384 285456 6390
rect 285404 6326 285456 6332
rect 284944 3120 284996 3126
rect 284944 3062 284996 3068
rect 285416 480 285444 6326
rect 286336 3398 286364 296210
rect 287072 9518 287100 301838
rect 287796 298716 287848 298722
rect 287796 298658 287848 298664
rect 287704 296540 287756 296546
rect 287704 296482 287756 296488
rect 287060 9512 287112 9518
rect 287060 9454 287112 9460
rect 286324 3392 286376 3398
rect 286324 3334 286376 3340
rect 286600 3392 286652 3398
rect 286600 3334 286652 3340
rect 286612 480 286640 3334
rect 287716 3330 287744 296482
rect 287808 11014 287836 298658
rect 288452 11830 288480 301838
rect 288728 299282 288756 301838
rect 288544 299254 288756 299282
rect 288544 49026 288572 299254
rect 288624 298376 288676 298382
rect 288624 298318 288676 298324
rect 288636 296614 288664 298318
rect 288624 296608 288676 296614
rect 288624 296550 288676 296556
rect 288532 49020 288584 49026
rect 288532 48962 288584 48968
rect 289084 14680 289136 14686
rect 289084 14622 289136 14628
rect 288440 11824 288492 11830
rect 288440 11766 288492 11772
rect 287796 11008 287848 11014
rect 287796 10950 287848 10956
rect 288992 6452 289044 6458
rect 288992 6394 289044 6400
rect 287704 3324 287756 3330
rect 287704 3266 287756 3272
rect 287796 3120 287848 3126
rect 287796 3062 287848 3068
rect 287808 480 287836 3062
rect 289004 480 289032 6394
rect 289096 3942 289124 14622
rect 289924 9654 289952 301838
rect 291028 298382 291056 301852
rect 291212 301838 291870 301866
rect 291016 298376 291068 298382
rect 291016 298318 291068 298324
rect 289912 9648 289964 9654
rect 289912 9590 289964 9596
rect 291212 7342 291240 301838
rect 291844 295928 291896 295934
rect 291844 295870 291896 295876
rect 291200 7336 291252 7342
rect 291200 7278 291252 7284
rect 291856 4010 291884 295870
rect 292684 8906 292712 301852
rect 293512 299470 293540 301852
rect 293972 301838 294354 301866
rect 294432 301838 295182 301866
rect 293500 299464 293552 299470
rect 293500 299406 293552 299412
rect 292672 8900 292724 8906
rect 292672 8842 292724 8848
rect 293972 6866 294000 301838
rect 294432 296714 294460 301838
rect 295904 299130 295932 301852
rect 296076 299464 296128 299470
rect 296076 299406 296128 299412
rect 295892 299124 295944 299130
rect 295892 299066 295944 299072
rect 295984 299124 296036 299130
rect 295984 299066 296036 299072
rect 294064 296686 294460 296714
rect 294064 7274 294092 296686
rect 294052 7268 294104 7274
rect 294052 7210 294104 7216
rect 293960 6860 294012 6866
rect 293960 6802 294012 6808
rect 292580 6520 292632 6526
rect 292580 6462 292632 6468
rect 291844 4004 291896 4010
rect 291844 3946 291896 3952
rect 289084 3936 289136 3942
rect 289084 3878 289136 3884
rect 290188 3324 290240 3330
rect 290188 3266 290240 3272
rect 290200 480 290228 3266
rect 291384 3256 291436 3262
rect 291384 3198 291436 3204
rect 291396 480 291424 3198
rect 292592 480 292620 6462
rect 293684 4004 293736 4010
rect 293684 3946 293736 3952
rect 293696 480 293724 3946
rect 294880 3188 294932 3194
rect 294880 3130 294932 3136
rect 294892 480 294920 3130
rect 295996 3126 296024 299066
rect 296088 10810 296116 299406
rect 296076 10804 296128 10810
rect 296076 10746 296128 10752
rect 296628 10532 296680 10538
rect 296628 10474 296680 10480
rect 295984 3120 296036 3126
rect 295984 3062 296036 3068
rect 296640 3058 296668 10474
rect 296732 6118 296760 301852
rect 296824 301838 297574 301866
rect 296824 7206 296852 301838
rect 298388 299334 298416 301852
rect 298572 301838 299230 301866
rect 299584 301838 300058 301866
rect 298376 299328 298428 299334
rect 298376 299270 298428 299276
rect 298572 296714 298600 301838
rect 298836 298648 298888 298654
rect 298836 298590 298888 298596
rect 298204 296686 298600 296714
rect 296812 7200 296864 7206
rect 296812 7142 296864 7148
rect 296720 6112 296772 6118
rect 296720 6054 296772 6060
rect 298204 6050 298232 296686
rect 298744 296336 298796 296342
rect 298744 296278 298796 296284
rect 298192 6044 298244 6050
rect 298192 5986 298244 5992
rect 298468 4072 298520 4078
rect 298468 4014 298520 4020
rect 297272 3256 297324 3262
rect 297272 3198 297324 3204
rect 296076 3052 296128 3058
rect 296076 2994 296128 3000
rect 296628 3052 296680 3058
rect 296628 2994 296680 3000
rect 296088 480 296116 2994
rect 297284 480 297312 3198
rect 298480 480 298508 4014
rect 298756 4010 298784 296278
rect 298848 10742 298876 298590
rect 298836 10736 298888 10742
rect 298836 10678 298888 10684
rect 299584 7138 299612 301838
rect 300124 299328 300176 299334
rect 300124 299270 300176 299276
rect 300136 12102 300164 299270
rect 300780 299198 300808 301852
rect 300872 301838 301622 301866
rect 302252 301838 302450 301866
rect 302712 301838 303278 301866
rect 303632 301838 304106 301866
rect 304184 301838 304842 301866
rect 305288 301838 305670 301866
rect 306392 301838 306498 301866
rect 306760 301838 307326 301866
rect 300768 299192 300820 299198
rect 300768 299134 300820 299140
rect 300124 12096 300176 12102
rect 300124 12038 300176 12044
rect 300768 11756 300820 11762
rect 300768 11698 300820 11704
rect 299572 7132 299624 7138
rect 299572 7074 299624 7080
rect 299664 5364 299716 5370
rect 299664 5306 299716 5312
rect 298744 4004 298796 4010
rect 298744 3946 298796 3952
rect 299676 480 299704 5306
rect 300780 480 300808 11698
rect 300872 5982 300900 301838
rect 302252 7070 302280 301838
rect 302712 296714 302740 301838
rect 302344 296686 302740 296714
rect 302344 11898 302372 296686
rect 302332 11892 302384 11898
rect 302332 11834 302384 11840
rect 302240 7064 302292 7070
rect 302240 7006 302292 7012
rect 300860 5976 300912 5982
rect 300860 5918 300912 5924
rect 303632 5914 303660 301838
rect 304184 299282 304212 301838
rect 303724 299254 304212 299282
rect 303724 296682 303752 299254
rect 305288 297362 305316 301838
rect 305828 298648 305880 298654
rect 305828 298590 305880 298596
rect 305644 298580 305696 298586
rect 305644 298522 305696 298528
rect 305276 297356 305328 297362
rect 305276 297298 305328 297304
rect 303712 296676 303764 296682
rect 303712 296618 303764 296624
rect 304264 296472 304316 296478
rect 304264 296414 304316 296420
rect 303620 5908 303672 5914
rect 303620 5850 303672 5856
rect 303160 5432 303212 5438
rect 303160 5374 303212 5380
rect 301964 3120 302016 3126
rect 301964 3062 302016 3068
rect 301976 480 302004 3062
rect 303172 480 303200 5374
rect 304276 3262 304304 296414
rect 305656 6914 305684 298522
rect 305736 297900 305788 297906
rect 305736 297842 305788 297848
rect 305472 6886 305684 6914
rect 305472 4146 305500 6886
rect 305460 4140 305512 4146
rect 305460 4082 305512 4088
rect 305552 4004 305604 4010
rect 305552 3946 305604 3952
rect 304264 3256 304316 3262
rect 304264 3198 304316 3204
rect 304356 3256 304408 3262
rect 304356 3198 304408 3204
rect 304368 480 304396 3198
rect 305564 480 305592 3946
rect 305748 3262 305776 297842
rect 305840 10674 305868 298590
rect 305828 10668 305880 10674
rect 305828 10610 305880 10616
rect 306392 5846 306420 301838
rect 306760 296714 306788 301838
rect 308140 299334 308168 301852
rect 308324 301838 308982 301866
rect 309152 301838 309718 301866
rect 308128 299328 308180 299334
rect 308128 299270 308180 299276
rect 308324 296714 308352 301838
rect 306484 296686 306788 296714
rect 307864 296686 308352 296714
rect 306484 11966 306512 296686
rect 306472 11960 306524 11966
rect 306472 11902 306524 11908
rect 306380 5840 306432 5846
rect 306380 5782 306432 5788
rect 307864 5778 307892 296686
rect 307852 5772 307904 5778
rect 307852 5714 307904 5720
rect 306748 5500 306800 5506
rect 306748 5442 306800 5448
rect 305736 3256 305788 3262
rect 305736 3198 305788 3204
rect 306760 480 306788 5442
rect 309152 4826 309180 301838
rect 310532 298654 310560 301852
rect 310624 301838 311374 301866
rect 310520 298648 310572 298654
rect 310520 298590 310572 298596
rect 309784 296676 309836 296682
rect 309784 296618 309836 296624
rect 309140 4820 309192 4826
rect 309140 4762 309192 4768
rect 309796 3330 309824 296618
rect 310624 6186 310652 301838
rect 312188 299198 312216 301852
rect 313016 299470 313044 301852
rect 313384 301838 313766 301866
rect 314304 301838 314594 301866
rect 313004 299464 313056 299470
rect 313004 299406 313056 299412
rect 313280 299328 313332 299334
rect 313280 299270 313332 299276
rect 312176 299192 312228 299198
rect 312176 299134 312228 299140
rect 312544 299192 312596 299198
rect 312544 299134 312596 299140
rect 312556 13122 312584 299134
rect 312636 18624 312688 18630
rect 312636 18566 312688 18572
rect 312544 13116 312596 13122
rect 312544 13058 312596 13064
rect 310612 6180 310664 6186
rect 310612 6122 310664 6128
rect 311624 6180 311676 6186
rect 311624 6122 311676 6128
rect 310244 4820 310296 4826
rect 310244 4762 310296 4768
rect 309784 3324 309836 3330
rect 309784 3266 309836 3272
rect 307944 3120 307996 3126
rect 307944 3062 307996 3068
rect 307956 480 307984 3062
rect 309048 2984 309100 2990
rect 309048 2926 309100 2932
rect 309060 480 309088 2926
rect 310256 480 310284 4762
rect 311440 3324 311492 3330
rect 311440 3266 311492 3272
rect 311452 480 311480 3266
rect 311636 3126 311664 6122
rect 312648 3330 312676 18566
rect 313292 4894 313320 299270
rect 313384 6254 313412 301838
rect 314304 299334 314332 301838
rect 314292 299328 314344 299334
rect 314292 299270 314344 299276
rect 315408 298722 315436 301852
rect 316052 301838 316250 301866
rect 316512 301838 317078 301866
rect 315396 298716 315448 298722
rect 315396 298658 315448 298664
rect 313372 6248 313424 6254
rect 313372 6190 313424 6196
rect 316052 5710 316080 301838
rect 316512 296714 316540 301838
rect 317892 299402 317920 301852
rect 317984 301838 318642 301866
rect 317880 299396 317932 299402
rect 317880 299338 317932 299344
rect 317420 298444 317472 298450
rect 317420 298386 317472 298392
rect 316144 296686 316540 296714
rect 316144 17270 316172 296686
rect 317432 294642 317460 298386
rect 317984 296714 318012 301838
rect 319456 299198 319484 301852
rect 320180 299328 320232 299334
rect 320180 299270 320232 299276
rect 319444 299192 319496 299198
rect 319444 299134 319496 299140
rect 317524 296686 318012 296714
rect 317420 294636 317472 294642
rect 317420 294578 317472 294584
rect 316132 17264 316184 17270
rect 316132 17206 316184 17212
rect 316040 5704 316092 5710
rect 316040 5646 316092 5652
rect 317524 5642 317552 296686
rect 318064 296608 318116 296614
rect 318064 296550 318116 296556
rect 317512 5636 317564 5642
rect 317512 5578 317564 5584
rect 313280 4888 313332 4894
rect 313280 4830 313332 4836
rect 313832 4888 313884 4894
rect 313832 4830 313884 4836
rect 312636 3324 312688 3330
rect 312636 3266 312688 3272
rect 312728 3324 312780 3330
rect 312728 3266 312780 3272
rect 311624 3120 311676 3126
rect 311624 3062 311676 3068
rect 312740 1714 312768 3266
rect 312648 1686 312768 1714
rect 312648 480 312676 1686
rect 313844 480 313872 4830
rect 317328 4752 317380 4758
rect 317328 4694 317380 4700
rect 316224 3256 316276 3262
rect 316224 3198 316276 3204
rect 315028 2916 315080 2922
rect 315028 2858 315080 2864
rect 315040 480 315068 2858
rect 316236 480 316264 3198
rect 317340 480 317368 4694
rect 318076 2922 318104 296550
rect 320192 5098 320220 299270
rect 320284 140078 320312 301852
rect 320744 301838 321126 301866
rect 321572 301838 321954 301866
rect 320744 299334 320772 301838
rect 320732 299328 320784 299334
rect 320732 299270 320784 299276
rect 320824 297356 320876 297362
rect 320824 297298 320876 297304
rect 320272 140072 320324 140078
rect 320272 140014 320324 140020
rect 320180 5092 320232 5098
rect 320180 5034 320232 5040
rect 319720 4140 319772 4146
rect 319720 4082 319772 4088
rect 318524 3052 318576 3058
rect 318524 2994 318576 3000
rect 318064 2916 318116 2922
rect 318064 2858 318116 2864
rect 318536 480 318564 2994
rect 319732 480 319760 4082
rect 320836 3398 320864 297298
rect 320916 5092 320968 5098
rect 320916 5034 320968 5040
rect 320824 3392 320876 3398
rect 320824 3334 320876 3340
rect 320928 480 320956 5034
rect 321572 4962 321600 301838
rect 322204 299192 322256 299198
rect 322204 299134 322256 299140
rect 321560 4956 321612 4962
rect 321560 4898 321612 4904
rect 322112 3392 322164 3398
rect 322112 3334 322164 3340
rect 322124 480 322152 3334
rect 322216 3262 322244 299134
rect 322676 297090 322704 301852
rect 322952 301838 323518 301866
rect 322664 297084 322716 297090
rect 322664 297026 322716 297032
rect 322952 5030 322980 301838
rect 323584 297968 323636 297974
rect 323584 297910 323636 297916
rect 322940 5024 322992 5030
rect 322940 4966 322992 4972
rect 323596 3398 323624 297910
rect 324332 8838 324360 301852
rect 324964 298648 325016 298654
rect 324964 298590 325016 298596
rect 324320 8832 324372 8838
rect 324320 8774 324372 8780
rect 324412 5024 324464 5030
rect 324412 4966 324464 4972
rect 323584 3392 323636 3398
rect 323584 3334 323636 3340
rect 322204 3256 322256 3262
rect 322204 3198 322256 3204
rect 323308 3256 323360 3262
rect 323308 3198 323360 3204
rect 323320 480 323348 3198
rect 324424 480 324452 4966
rect 324976 3126 325004 298590
rect 325160 297022 325188 301852
rect 325804 301838 326002 301866
rect 326448 301838 326830 301866
rect 325700 299328 325752 299334
rect 325700 299270 325752 299276
rect 325148 297016 325200 297022
rect 325148 296958 325200 296964
rect 325712 8702 325740 299270
rect 325804 296002 325832 301838
rect 326448 299334 326476 301838
rect 326436 299328 326488 299334
rect 326436 299270 326488 299276
rect 327552 296954 327580 301852
rect 327644 301838 328394 301866
rect 328472 301838 329222 301866
rect 327540 296948 327592 296954
rect 327540 296890 327592 296896
rect 327644 296714 327672 301838
rect 327724 299328 327776 299334
rect 327724 299270 327776 299276
rect 327092 296686 327672 296714
rect 325792 295996 325844 296002
rect 325792 295938 325844 295944
rect 325700 8696 325752 8702
rect 325700 8638 325752 8644
rect 327092 5166 327120 296686
rect 327080 5160 327132 5166
rect 327080 5102 327132 5108
rect 326804 3324 326856 3330
rect 326804 3266 326856 3272
rect 324964 3120 325016 3126
rect 324964 3062 325016 3068
rect 325608 3120 325660 3126
rect 325608 3062 325660 3068
rect 325620 480 325648 3062
rect 326816 480 326844 3266
rect 327736 3262 327764 299270
rect 328472 8770 328500 301838
rect 329104 298716 329156 298722
rect 329104 298658 329156 298664
rect 328460 8764 328512 8770
rect 328460 8706 328512 8712
rect 328000 4956 328052 4962
rect 328000 4898 328052 4904
rect 327724 3256 327776 3262
rect 327724 3198 327776 3204
rect 328012 480 328040 4898
rect 329116 2990 329144 298658
rect 330036 298042 330064 301852
rect 330312 301838 330878 301866
rect 331232 301838 331614 301866
rect 330024 298036 330076 298042
rect 330024 297978 330076 297984
rect 330312 296714 330340 301838
rect 329852 296686 330340 296714
rect 329852 5234 329880 296686
rect 331232 8634 331260 301838
rect 331864 299396 331916 299402
rect 331864 299338 331916 299344
rect 331220 8628 331272 8634
rect 331220 8570 331272 8576
rect 329840 5228 329892 5234
rect 329840 5170 329892 5176
rect 331588 5160 331640 5166
rect 331588 5102 331640 5108
rect 330392 3392 330444 3398
rect 330392 3334 330444 3340
rect 329104 2984 329156 2990
rect 329104 2926 329156 2932
rect 329196 2916 329248 2922
rect 329196 2858 329248 2864
rect 329208 480 329236 2858
rect 330404 480 330432 3334
rect 331600 480 331628 5102
rect 331876 3398 331904 299338
rect 332428 297158 332456 301852
rect 332612 301838 333270 301866
rect 333992 301838 334098 301866
rect 334452 301838 334926 301866
rect 335464 301838 335754 301866
rect 336200 301838 336490 301866
rect 332416 297152 332468 297158
rect 332416 297094 332468 297100
rect 332612 295798 332640 301838
rect 332600 295792 332652 295798
rect 332600 295734 332652 295740
rect 333992 8566 334020 301838
rect 334452 296714 334480 301838
rect 335360 299464 335412 299470
rect 335360 299406 335412 299412
rect 334084 296686 334480 296714
rect 334084 13190 334112 296686
rect 334072 13184 334124 13190
rect 334072 13126 334124 13132
rect 333980 8560 334032 8566
rect 333980 8502 334032 8508
rect 335372 8430 335400 299406
rect 335464 296070 335492 301838
rect 336200 299470 336228 301838
rect 336188 299464 336240 299470
rect 336188 299406 336240 299412
rect 337304 297226 337332 301852
rect 338146 301838 338252 301866
rect 338120 299464 338172 299470
rect 338120 299406 338172 299412
rect 338028 298376 338080 298382
rect 338028 298318 338080 298324
rect 337292 297220 337344 297226
rect 337292 297162 337344 297168
rect 335452 296064 335504 296070
rect 335452 296006 335504 296012
rect 336648 295996 336700 296002
rect 336648 295938 336700 295944
rect 335360 8424 335412 8430
rect 335360 8366 335412 8372
rect 335084 5228 335136 5234
rect 335084 5170 335136 5176
rect 331864 3392 331916 3398
rect 331864 3334 331916 3340
rect 332692 2984 332744 2990
rect 332692 2926 332744 2932
rect 332704 480 332732 2926
rect 333888 2848 333940 2854
rect 333888 2790 333940 2796
rect 333900 480 333928 2790
rect 335096 480 335124 5170
rect 336292 598 336504 626
rect 336292 480 336320 598
rect 336476 490 336504 598
rect 336660 490 336688 295938
rect 338040 6914 338068 298318
rect 338132 8498 338160 299406
rect 338224 295866 338252 301838
rect 338592 301838 338974 301866
rect 339604 301838 339802 301866
rect 340248 301838 340538 301866
rect 338592 299470 338620 301838
rect 338580 299464 338632 299470
rect 338580 299406 338632 299412
rect 339500 299464 339552 299470
rect 339500 299406 339552 299412
rect 338764 298512 338816 298518
rect 338764 298454 338816 298460
rect 338212 295860 338264 295866
rect 338212 295802 338264 295808
rect 338120 8492 338172 8498
rect 338120 8434 338172 8440
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 336476 462 336688 490
rect 337488 6886 338068 6914
rect 337488 480 337516 6886
rect 338672 4684 338724 4690
rect 338672 4626 338724 4632
rect 338684 480 338712 4626
rect 338776 3194 338804 298454
rect 339512 5302 339540 299406
rect 339604 14482 339632 301838
rect 340248 299470 340276 301838
rect 340236 299464 340288 299470
rect 340236 299406 340288 299412
rect 341352 298450 341380 301852
rect 341444 301838 342194 301866
rect 342272 301838 343022 301866
rect 343652 301838 343850 301866
rect 341340 298444 341392 298450
rect 341340 298386 341392 298392
rect 341444 296714 341472 301838
rect 341524 298104 341576 298110
rect 341524 298046 341576 298052
rect 340984 296686 341472 296714
rect 340984 141438 341012 296686
rect 340972 141432 341024 141438
rect 340972 141374 341024 141380
rect 339592 14476 339644 14482
rect 339592 14418 339644 14424
rect 339868 6588 339920 6594
rect 339868 6530 339920 6536
rect 339500 5296 339552 5302
rect 339500 5238 339552 5244
rect 338764 3188 338816 3194
rect 338764 3130 338816 3136
rect 339880 480 339908 6530
rect 340972 3188 341024 3194
rect 340972 3130 341024 3136
rect 340984 480 341012 3130
rect 341536 2854 341564 298046
rect 342272 7682 342300 301838
rect 343548 298036 343600 298042
rect 343548 297978 343600 297984
rect 342260 7676 342312 7682
rect 342260 7618 342312 7624
rect 343560 6914 343588 297978
rect 343652 296138 343680 301838
rect 344664 297430 344692 301852
rect 345124 301838 345414 301866
rect 344652 297424 344704 297430
rect 344652 297366 344704 297372
rect 343640 296132 343692 296138
rect 343640 296074 343692 296080
rect 345124 7614 345152 301838
rect 346228 298858 346256 301852
rect 346688 301838 347070 301866
rect 346216 298852 346268 298858
rect 346216 298794 346268 298800
rect 345664 298444 345716 298450
rect 345664 298386 345716 298392
rect 345112 7608 345164 7614
rect 345112 7550 345164 7556
rect 343376 6886 343588 6914
rect 342168 5296 342220 5302
rect 342168 5238 342220 5244
rect 341524 2848 341576 2854
rect 341524 2790 341576 2796
rect 342180 480 342208 5238
rect 343376 480 343404 6886
rect 345676 3466 345704 298386
rect 346688 297498 346716 301838
rect 347044 298920 347096 298926
rect 347044 298862 347096 298868
rect 346676 297492 346728 297498
rect 346676 297434 346728 297440
rect 346952 6248 347004 6254
rect 346952 6190 347004 6196
rect 345756 4616 345808 4622
rect 345756 4558 345808 4564
rect 344560 3460 344612 3466
rect 344560 3402 344612 3408
rect 345664 3460 345716 3466
rect 345664 3402 345716 3408
rect 344572 480 344600 3402
rect 345768 480 345796 4558
rect 346964 480 346992 6190
rect 347056 2922 347084 298862
rect 347884 7750 347912 301852
rect 348712 298926 348740 301852
rect 348700 298920 348752 298926
rect 348700 298862 348752 298868
rect 349448 297838 349476 301852
rect 349540 301838 350290 301866
rect 349436 297832 349488 297838
rect 349436 297774 349488 297780
rect 349540 296714 349568 301838
rect 351104 298858 351132 301852
rect 351946 301838 352052 301866
rect 351920 299532 351972 299538
rect 351920 299474 351972 299480
rect 351828 298920 351880 298926
rect 351828 298862 351880 298868
rect 351092 298852 351144 298858
rect 351092 298794 351144 298800
rect 350356 297424 350408 297430
rect 350356 297366 350408 297372
rect 349172 296686 349568 296714
rect 349172 7818 349200 296686
rect 350368 16574 350396 297366
rect 350368 16546 350488 16574
rect 349160 7812 349212 7818
rect 349160 7754 349212 7760
rect 347872 7744 347924 7750
rect 347872 7686 347924 7692
rect 349252 4548 349304 4554
rect 349252 4490 349304 4496
rect 348056 3460 348108 3466
rect 348056 3402 348108 3408
rect 347044 2916 347096 2922
rect 347044 2858 347096 2864
rect 348068 480 348096 3402
rect 349264 480 349292 4490
rect 350460 480 350488 16546
rect 351840 6914 351868 298862
rect 351932 7886 351960 299474
rect 352024 10606 352052 301838
rect 352392 301838 352774 301866
rect 353496 301838 353602 301866
rect 354048 301838 354338 301866
rect 354784 301838 355166 301866
rect 352392 299538 352420 301838
rect 352380 299532 352432 299538
rect 352380 299474 352432 299480
rect 353392 299532 353444 299538
rect 353392 299474 353444 299480
rect 353404 12170 353432 299474
rect 353392 12164 353444 12170
rect 353392 12106 353444 12112
rect 352012 10600 352064 10606
rect 352012 10542 352064 10548
rect 351920 7880 351972 7886
rect 351920 7822 351972 7828
rect 351656 6886 351868 6914
rect 351656 480 351684 6886
rect 352840 4480 352892 4486
rect 352840 4422 352892 4428
rect 352852 480 352880 4422
rect 353496 3534 353524 301838
rect 354048 299538 354076 301838
rect 354036 299532 354088 299538
rect 354036 299474 354088 299480
rect 354588 11824 354640 11830
rect 354588 11766 354640 11772
rect 354600 3534 354628 11766
rect 354784 7954 354812 301838
rect 355980 299266 356008 301852
rect 356072 301838 356822 301866
rect 357544 301838 357650 301866
rect 358096 301838 358478 301866
rect 358924 301838 359214 301866
rect 359752 301838 360042 301866
rect 355968 299260 356020 299266
rect 355968 299202 356020 299208
rect 356072 10878 356100 301838
rect 357440 299260 357492 299266
rect 357440 299202 357492 299208
rect 356704 297288 356756 297294
rect 356704 297230 356756 297236
rect 356060 10872 356112 10878
rect 356060 10814 356112 10820
rect 354772 7948 354824 7954
rect 354772 7890 354824 7896
rect 356336 4412 356388 4418
rect 356336 4354 356388 4360
rect 355232 3664 355284 3670
rect 355232 3606 355284 3612
rect 353484 3528 353536 3534
rect 353484 3470 353536 3476
rect 354036 3528 354088 3534
rect 354036 3470 354088 3476
rect 354588 3528 354640 3534
rect 354588 3470 354640 3476
rect 354048 480 354076 3470
rect 355244 480 355272 3606
rect 356348 480 356376 4354
rect 356716 2990 356744 297230
rect 357452 3602 357480 299202
rect 357544 296410 357572 301838
rect 358096 299266 358124 301838
rect 358084 299260 358136 299266
rect 358084 299202 358136 299208
rect 358820 299260 358872 299266
rect 358820 299202 358872 299208
rect 358728 298444 358780 298450
rect 358728 298386 358780 298392
rect 357532 296404 357584 296410
rect 357532 296346 357584 296352
rect 357440 3596 357492 3602
rect 357440 3538 357492 3544
rect 356704 2984 356756 2990
rect 356704 2926 356756 2932
rect 357532 2984 357584 2990
rect 357532 2926 357584 2932
rect 357544 480 357572 2926
rect 358740 480 358768 298386
rect 358832 10946 358860 299202
rect 358924 14618 358952 301838
rect 359752 299266 359780 301838
rect 359740 299260 359792 299266
rect 359740 299202 359792 299208
rect 360856 298586 360884 301852
rect 360844 298580 360896 298586
rect 360844 298522 360896 298528
rect 360844 297832 360896 297838
rect 360844 297774 360896 297780
rect 358912 14612 358964 14618
rect 358912 14554 358964 14560
rect 359464 11892 359516 11898
rect 359464 11834 359516 11840
rect 358820 10940 358872 10946
rect 358820 10882 358872 10888
rect 359476 2990 359504 11834
rect 359924 4344 359976 4350
rect 359924 4286 359976 4292
rect 359464 2984 359516 2990
rect 359464 2926 359516 2932
rect 359936 480 359964 4286
rect 360856 3058 360884 297774
rect 361684 297702 361712 301852
rect 361960 301838 362526 301866
rect 361672 297696 361724 297702
rect 361672 297638 361724 297644
rect 361960 296714 361988 301838
rect 363248 299266 363276 301852
rect 363524 301838 364090 301866
rect 364352 301838 364918 301866
rect 362224 299260 362276 299266
rect 362224 299202 362276 299208
rect 363236 299260 363288 299266
rect 363236 299202 363288 299208
rect 361592 296686 361988 296714
rect 361592 296206 361620 296686
rect 361580 296200 361632 296206
rect 361580 296142 361632 296148
rect 362236 3602 362264 299202
rect 363524 296714 363552 301838
rect 363064 296686 363552 296714
rect 363064 10402 363092 296686
rect 364352 14550 364380 301838
rect 365732 298790 365760 301852
rect 365720 298784 365772 298790
rect 365720 298726 365772 298732
rect 366560 297634 366588 301852
rect 367204 301838 367402 301866
rect 367848 301838 368138 301866
rect 367100 299532 367152 299538
rect 367100 299474 367152 299480
rect 366548 297628 366600 297634
rect 366548 297570 366600 297576
rect 364340 14544 364392 14550
rect 364340 14486 364392 14492
rect 363052 10396 363104 10402
rect 363052 10338 363104 10344
rect 363604 10396 363656 10402
rect 363604 10338 363656 10344
rect 363512 4276 363564 4282
rect 363512 4218 363564 4224
rect 362224 3596 362276 3602
rect 362224 3538 362276 3544
rect 362316 3596 362368 3602
rect 362316 3538 362368 3544
rect 361120 3528 361172 3534
rect 361120 3470 361172 3476
rect 360844 3052 360896 3058
rect 360844 2994 360896 3000
rect 361132 480 361160 3470
rect 362328 480 362356 3538
rect 363524 480 363552 4218
rect 363616 3534 363644 10338
rect 367008 6656 367060 6662
rect 367008 6598 367060 6604
rect 365812 3664 365864 3670
rect 365812 3606 365864 3612
rect 363604 3528 363656 3534
rect 363604 3470 363656 3476
rect 364616 2984 364668 2990
rect 364616 2926 364668 2932
rect 364628 480 364656 2926
rect 365824 480 365852 3606
rect 367020 480 367048 6598
rect 367112 3738 367140 299474
rect 367204 202162 367232 301838
rect 367848 299538 367876 301838
rect 367836 299532 367888 299538
rect 367836 299474 367888 299480
rect 367744 298784 367796 298790
rect 367744 298726 367796 298732
rect 367192 202156 367244 202162
rect 367192 202098 367244 202104
rect 367100 3732 367152 3738
rect 367100 3674 367152 3680
rect 367756 3670 367784 298726
rect 368952 297566 368980 301852
rect 369136 301838 369794 301866
rect 368940 297560 368992 297566
rect 368940 297502 368992 297508
rect 369136 296714 369164 301838
rect 370608 299062 370636 301852
rect 371252 301838 371450 301866
rect 371804 301838 372186 301866
rect 370596 299056 370648 299062
rect 370596 298998 370648 299004
rect 370504 297220 370556 297226
rect 370504 297162 370556 297168
rect 368492 296686 369164 296714
rect 368492 296546 368520 296686
rect 368480 296540 368532 296546
rect 368480 296482 368532 296488
rect 369400 3732 369452 3738
rect 369400 3674 369452 3680
rect 367744 3664 367796 3670
rect 367744 3606 367796 3612
rect 368204 3664 368256 3670
rect 368204 3606 368256 3612
rect 368216 480 368244 3606
rect 369412 480 369440 3674
rect 370516 3126 370544 297162
rect 370596 296132 370648 296138
rect 370596 296074 370648 296080
rect 370608 3670 370636 296074
rect 371252 10470 371280 301838
rect 371804 296714 371832 301838
rect 373000 299062 373028 301852
rect 371884 299056 371936 299062
rect 371884 298998 371936 299004
rect 372988 299056 373040 299062
rect 372988 298998 373040 299004
rect 371344 296686 371832 296714
rect 371344 295934 371372 296686
rect 371332 295928 371384 295934
rect 371332 295870 371384 295876
rect 371240 10464 371292 10470
rect 371240 10406 371292 10412
rect 371700 7608 371752 7614
rect 371700 7550 371752 7556
rect 370688 6724 370740 6730
rect 370688 6666 370740 6672
rect 370596 3664 370648 3670
rect 370596 3606 370648 3612
rect 370700 3210 370728 6666
rect 370608 3182 370728 3210
rect 370504 3120 370556 3126
rect 370504 3062 370556 3068
rect 370608 480 370636 3182
rect 371712 480 371740 7550
rect 371896 3806 371924 298998
rect 373828 297770 373856 301852
rect 374012 301838 374670 301866
rect 373908 299056 373960 299062
rect 373908 298998 373960 299004
rect 373816 297764 373868 297770
rect 373816 297706 373868 297712
rect 371884 3800 371936 3806
rect 371884 3742 371936 3748
rect 373920 3738 373948 298998
rect 374012 14686 374040 301838
rect 375484 298994 375512 301852
rect 375760 301838 376326 301866
rect 376864 301838 377062 301866
rect 377600 301838 377890 301866
rect 378152 301838 378718 301866
rect 375472 298988 375524 298994
rect 375472 298930 375524 298936
rect 375760 296714 375788 301838
rect 376760 299124 376812 299130
rect 376760 299066 376812 299072
rect 375484 296686 375788 296714
rect 375288 296064 375340 296070
rect 375288 296006 375340 296012
rect 374000 14680 374052 14686
rect 374000 14622 374052 14628
rect 374092 6792 374144 6798
rect 374092 6734 374144 6740
rect 372896 3732 372948 3738
rect 372896 3674 372948 3680
rect 373908 3732 373960 3738
rect 373908 3674 373960 3680
rect 372908 480 372936 3674
rect 374104 480 374132 6734
rect 375300 480 375328 296006
rect 375484 6322 375512 296686
rect 376024 296200 376076 296206
rect 376024 296142 376076 296148
rect 375472 6316 375524 6322
rect 375472 6258 375524 6264
rect 376036 2990 376064 296142
rect 376772 3874 376800 299066
rect 376864 296274 376892 301838
rect 377600 299130 377628 301838
rect 377588 299124 377640 299130
rect 377588 299066 377640 299072
rect 378048 297492 378100 297498
rect 378048 297434 378100 297440
rect 376852 296268 376904 296274
rect 376852 296210 376904 296216
rect 376760 3868 376812 3874
rect 376760 3810 376812 3816
rect 376484 3120 376536 3126
rect 376484 3062 376536 3068
rect 376024 2984 376076 2990
rect 376024 2926 376076 2932
rect 376496 480 376524 3062
rect 377692 598 377904 626
rect 377692 480 377720 598
rect 377876 490 377904 598
rect 378060 490 378088 297434
rect 378152 6390 378180 301838
rect 379532 297362 379560 301852
rect 380164 299124 380216 299130
rect 380164 299066 380216 299072
rect 379520 297356 379572 297362
rect 379520 297298 379572 297304
rect 378140 6384 378192 6390
rect 378140 6326 378192 6332
rect 380176 3806 380204 299066
rect 380360 298994 380388 301852
rect 380912 301838 381110 301866
rect 381188 301838 381938 301866
rect 382292 301838 382766 301866
rect 383304 301838 383594 301866
rect 383672 301838 384422 301866
rect 380348 298988 380400 298994
rect 380348 298930 380400 298936
rect 380808 298988 380860 298994
rect 380808 298930 380860 298936
rect 378876 3800 378928 3806
rect 378876 3742 378928 3748
rect 380164 3800 380216 3806
rect 380164 3742 380216 3748
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 377876 462 378088 490
rect 378888 480 378916 3742
rect 380820 3738 380848 298930
rect 380912 6458 380940 301838
rect 381188 299282 381216 301838
rect 381004 299254 381216 299282
rect 381004 296682 381032 299254
rect 382188 297560 382240 297566
rect 382188 297502 382240 297508
rect 380992 296676 381044 296682
rect 380992 296618 381044 296624
rect 380900 6452 380952 6458
rect 380900 6394 380952 6400
rect 382200 3738 382228 297502
rect 382292 3942 382320 301838
rect 383304 296714 383332 301838
rect 382384 296686 383332 296714
rect 382384 6526 382412 296686
rect 383672 296342 383700 301838
rect 384304 298648 384356 298654
rect 384304 298590 384356 298596
rect 383660 296336 383712 296342
rect 383660 296278 383712 296284
rect 382372 6520 382424 6526
rect 382372 6462 382424 6468
rect 382372 6384 382424 6390
rect 382372 6326 382424 6332
rect 382280 3936 382332 3942
rect 382280 3878 382332 3884
rect 379980 3732 380032 3738
rect 379980 3674 380032 3680
rect 380808 3732 380860 3738
rect 380808 3674 380860 3680
rect 381176 3732 381228 3738
rect 381176 3674 381228 3680
rect 382188 3732 382240 3738
rect 382188 3674 382240 3680
rect 379992 480 380020 3674
rect 381188 480 381216 3674
rect 382384 480 382412 6326
rect 384316 3874 384344 298590
rect 385236 298518 385264 301852
rect 385512 301838 385986 301866
rect 386524 301838 386814 301866
rect 385224 298512 385276 298518
rect 385224 298454 385276 298460
rect 385512 296714 385540 301838
rect 386328 298512 386380 298518
rect 386328 298454 386380 298460
rect 385144 296686 385540 296714
rect 385144 10538 385172 296686
rect 385132 10532 385184 10538
rect 385132 10474 385184 10480
rect 384764 6316 384816 6322
rect 384764 6258 384816 6264
rect 384304 3868 384356 3874
rect 384304 3810 384356 3816
rect 383568 3800 383620 3806
rect 383568 3742 383620 3748
rect 383580 480 383608 3742
rect 384776 480 384804 6258
rect 385972 598 386184 626
rect 385972 480 386000 598
rect 386156 490 386184 598
rect 386340 490 386368 298454
rect 386524 296478 386552 301838
rect 387628 298654 387656 301852
rect 387812 301838 388470 301866
rect 387616 298648 387668 298654
rect 387616 298590 387668 298596
rect 387708 298444 387760 298450
rect 387708 298386 387760 298392
rect 386512 296472 386564 296478
rect 386512 296414 386564 296420
rect 387720 3058 387748 298386
rect 387812 5370 387840 301838
rect 389284 11762 389312 301852
rect 390020 298586 390048 301852
rect 390572 301838 390862 301866
rect 390008 298580 390060 298586
rect 390008 298522 390060 298528
rect 389824 297628 389876 297634
rect 389824 297570 389876 297576
rect 389272 11756 389324 11762
rect 389272 11698 389324 11704
rect 389456 6452 389508 6458
rect 389456 6394 389508 6400
rect 387800 5364 387852 5370
rect 387800 5306 387852 5312
rect 387156 3052 387208 3058
rect 387156 2994 387208 3000
rect 387708 3052 387760 3058
rect 387708 2994 387760 3000
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386156 462 386368 490
rect 387168 480 387196 2994
rect 388260 2916 388312 2922
rect 388260 2858 388312 2864
rect 388272 480 388300 2858
rect 389468 480 389496 6394
rect 389836 2922 389864 297570
rect 390572 5438 390600 301838
rect 391204 298648 391256 298654
rect 391204 298590 391256 298596
rect 390560 5432 390612 5438
rect 390560 5374 390612 5380
rect 391216 4010 391244 298590
rect 391676 297906 391704 301852
rect 392504 298654 392532 301852
rect 392492 298648 392544 298654
rect 392492 298590 392544 298596
rect 392584 298648 392636 298654
rect 392584 298590 392636 298596
rect 391664 297900 391716 297906
rect 391664 297842 391716 297848
rect 391204 4004 391256 4010
rect 391204 3946 391256 3952
rect 392596 3942 392624 298590
rect 392676 297696 392728 297702
rect 392676 297638 392728 297644
rect 392584 3936 392636 3942
rect 392584 3878 392636 3884
rect 390652 3868 390704 3874
rect 390652 3810 390704 3816
rect 389824 2916 389876 2922
rect 389824 2858 389876 2864
rect 390664 480 390692 3810
rect 392688 3330 392716 297638
rect 393332 5506 393360 301852
rect 393424 301838 394174 301866
rect 393424 6186 393452 301838
rect 394896 298722 394924 301852
rect 395264 301838 395738 301866
rect 396184 301838 396566 301866
rect 394884 298716 394936 298722
rect 394884 298658 394936 298664
rect 395264 296714 395292 301838
rect 395988 297764 396040 297770
rect 395988 297706 396040 297712
rect 394804 296686 395292 296714
rect 393412 6180 393464 6186
rect 393412 6122 393464 6128
rect 393320 5500 393372 5506
rect 393320 5442 393372 5448
rect 394804 4826 394832 296686
rect 394792 4820 394844 4826
rect 394792 4762 394844 4768
rect 393044 4004 393096 4010
rect 393044 3946 393096 3952
rect 391848 3324 391900 3330
rect 391848 3266 391900 3272
rect 392676 3324 392728 3330
rect 392676 3266 392728 3272
rect 391860 480 391888 3266
rect 393056 480 393084 3946
rect 396000 3330 396028 297706
rect 396184 18630 396212 301838
rect 396724 298716 396776 298722
rect 396724 298658 396776 298664
rect 396172 18624 396224 18630
rect 396172 18566 396224 18572
rect 395344 3324 395396 3330
rect 395344 3266 395396 3272
rect 395988 3324 396040 3330
rect 395988 3266 396040 3272
rect 394240 3120 394292 3126
rect 394240 3062 394292 3068
rect 394252 480 394280 3062
rect 395356 480 395384 3266
rect 396736 3126 396764 298658
rect 397380 298654 397408 301852
rect 397472 301838 398222 301866
rect 397368 298648 397420 298654
rect 397368 298590 397420 298596
rect 396816 298512 396868 298518
rect 396816 298454 396868 298460
rect 396828 4010 396856 298454
rect 397472 4894 397500 301838
rect 398944 296614 398972 301852
rect 399404 301838 399786 301866
rect 400232 301838 400614 301866
rect 399404 299198 399432 301838
rect 399392 299192 399444 299198
rect 399392 299134 399444 299140
rect 399484 299192 399536 299198
rect 399484 299134 399536 299140
rect 398932 296608 398984 296614
rect 398932 296550 398984 296556
rect 397460 4888 397512 4894
rect 397460 4830 397512 4836
rect 399496 4146 399524 299134
rect 400128 298376 400180 298382
rect 400128 298318 400180 298324
rect 399484 4140 399536 4146
rect 399484 4082 399536 4088
rect 396816 4004 396868 4010
rect 396816 3946 396868 3952
rect 397736 4004 397788 4010
rect 397736 3946 397788 3952
rect 396724 3120 396776 3126
rect 396724 3062 396776 3068
rect 396540 3052 396592 3058
rect 396540 2994 396592 3000
rect 396552 480 396580 2994
rect 397748 480 397776 3946
rect 398932 3324 398984 3330
rect 398932 3266 398984 3272
rect 398944 480 398972 3266
rect 400140 480 400168 298318
rect 400232 4758 400260 301838
rect 401428 297906 401456 301852
rect 402256 299198 402284 301852
rect 402992 301838 403098 301866
rect 402244 299192 402296 299198
rect 402244 299134 402296 299140
rect 402244 298648 402296 298654
rect 402244 298590 402296 298596
rect 401416 297900 401468 297906
rect 401416 297842 401468 297848
rect 400864 297832 400916 297838
rect 400864 297774 400916 297780
rect 400220 4752 400272 4758
rect 400220 4694 400272 4700
rect 400876 3330 400904 297774
rect 402256 3330 402284 298590
rect 402992 5098 403020 301838
rect 403820 297974 403848 301852
rect 404648 299334 404676 301852
rect 404740 301838 405490 301866
rect 404636 299328 404688 299334
rect 404636 299270 404688 299276
rect 403808 297968 403860 297974
rect 403808 297910 403860 297916
rect 403624 297900 403676 297906
rect 403624 297842 403676 297848
rect 403636 6914 403664 297842
rect 404740 296714 404768 301838
rect 406304 297226 406332 301852
rect 407132 298246 407160 301852
rect 407224 301838 407882 301866
rect 406384 298240 406436 298246
rect 406384 298182 406436 298188
rect 407120 298240 407172 298246
rect 407120 298182 407172 298188
rect 406292 297220 406344 297226
rect 406292 297162 406344 297168
rect 403544 6886 403664 6914
rect 404464 296686 404768 296714
rect 402980 5092 403032 5098
rect 402980 5034 403032 5040
rect 403544 4146 403572 6886
rect 404464 5030 404492 296686
rect 404452 5024 404504 5030
rect 404452 4966 404504 4972
rect 402520 4140 402572 4146
rect 402520 4082 402572 4088
rect 403532 4140 403584 4146
rect 403532 4082 403584 4088
rect 400864 3324 400916 3330
rect 400864 3266 400916 3272
rect 401324 3324 401376 3330
rect 401324 3266 401376 3272
rect 402244 3324 402296 3330
rect 402244 3266 402296 3272
rect 401336 480 401364 3266
rect 402532 480 402560 4082
rect 403624 4072 403676 4078
rect 403624 4014 403676 4020
rect 403636 480 403664 4014
rect 406016 3392 406068 3398
rect 406016 3334 406068 3340
rect 404820 3324 404872 3330
rect 404820 3266 404872 3272
rect 404832 480 404860 3266
rect 406028 480 406056 3334
rect 406396 3262 406424 298182
rect 407028 297968 407080 297974
rect 407028 297910 407080 297916
rect 407040 3398 407068 297910
rect 407224 4962 407252 301838
rect 408408 299328 408460 299334
rect 408408 299270 408460 299276
rect 407212 4956 407264 4962
rect 407212 4898 407264 4904
rect 407028 3392 407080 3398
rect 407028 3334 407080 3340
rect 407212 3392 407264 3398
rect 407212 3334 407264 3340
rect 406384 3256 406436 3262
rect 406384 3198 406436 3204
rect 407224 480 407252 3334
rect 408420 480 408448 299270
rect 408696 298110 408724 301852
rect 409524 299402 409552 301852
rect 409892 301838 410366 301866
rect 409512 299396 409564 299402
rect 409512 299338 409564 299344
rect 408684 298104 408736 298110
rect 408684 298046 408736 298052
rect 409892 5166 409920 301838
rect 410524 299396 410576 299402
rect 410524 299338 410576 299344
rect 410536 6594 410564 299338
rect 411180 297294 411208 301852
rect 411272 301838 412022 301866
rect 412652 301838 412758 301866
rect 412836 301838 413586 301866
rect 411168 297288 411220 297294
rect 411168 297230 411220 297236
rect 410524 6588 410576 6594
rect 410524 6530 410576 6536
rect 409880 5160 409932 5166
rect 409880 5102 409932 5108
rect 410800 3256 410852 3262
rect 410800 3198 410852 3204
rect 409604 3052 409656 3058
rect 409604 2994 409656 3000
rect 409616 480 409644 2994
rect 410812 480 410840 3198
rect 411272 3126 411300 301838
rect 411904 298376 411956 298382
rect 411904 298318 411956 298324
rect 411916 3398 411944 298318
rect 412652 5234 412680 301838
rect 412836 296714 412864 301838
rect 414400 299470 414428 301852
rect 414492 301838 415242 301866
rect 414388 299464 414440 299470
rect 414388 299406 414440 299412
rect 413284 298104 413336 298110
rect 413284 298046 413336 298052
rect 412744 296686 412864 296714
rect 412744 296002 412772 296686
rect 412732 295996 412784 296002
rect 412732 295938 412784 295944
rect 412640 5228 412692 5234
rect 412640 5170 412692 5176
rect 413100 3460 413152 3466
rect 413100 3402 413152 3408
rect 411904 3392 411956 3398
rect 411904 3334 411956 3340
rect 411260 3120 411312 3126
rect 411260 3062 411312 3068
rect 411904 3120 411956 3126
rect 411904 3062 411956 3068
rect 411916 480 411944 3062
rect 413112 480 413140 3402
rect 413296 3058 413324 298046
rect 414492 296714 414520 301838
rect 416056 299402 416084 301852
rect 416792 301838 416898 301866
rect 417160 301838 417634 301866
rect 416688 299464 416740 299470
rect 416688 299406 416740 299412
rect 416044 299396 416096 299402
rect 416044 299338 416096 299344
rect 416044 298308 416096 298314
rect 416044 298250 416096 298256
rect 414664 297356 414716 297362
rect 414664 297298 414716 297304
rect 414124 296686 414520 296714
rect 414124 4690 414152 296686
rect 414112 4684 414164 4690
rect 414112 4626 414164 4632
rect 414676 3466 414704 297298
rect 414664 3460 414716 3466
rect 414664 3402 414716 3408
rect 415492 3460 415544 3466
rect 415492 3402 415544 3408
rect 414296 3392 414348 3398
rect 414296 3334 414348 3340
rect 413284 3052 413336 3058
rect 413284 2994 413336 3000
rect 414308 480 414336 3334
rect 415504 480 415532 3402
rect 416056 3398 416084 298250
rect 416700 3466 416728 299406
rect 416688 3460 416740 3466
rect 416688 3402 416740 3408
rect 416044 3392 416096 3398
rect 416044 3334 416096 3340
rect 416688 3256 416740 3262
rect 416688 3198 416740 3204
rect 416700 480 416728 3198
rect 416792 3194 416820 301838
rect 417160 296714 417188 301838
rect 418448 298042 418476 301852
rect 419276 298858 419304 301852
rect 419552 301838 420118 301866
rect 420946 301838 421052 301866
rect 419264 298852 419316 298858
rect 419264 298794 419316 298800
rect 418436 298036 418488 298042
rect 418436 297978 418488 297984
rect 418804 298036 418856 298042
rect 418804 297978 418856 297984
rect 416884 296686 417188 296714
rect 416884 5302 416912 296686
rect 416872 5296 416924 5302
rect 416872 5238 416924 5244
rect 418816 3262 418844 297978
rect 419552 4622 419580 301838
rect 420920 299396 420972 299402
rect 420920 299338 420972 299344
rect 420184 4820 420236 4826
rect 420184 4762 420236 4768
rect 419540 4616 419592 4622
rect 419540 4558 419592 4564
rect 418804 3256 418856 3262
rect 418804 3198 418856 3204
rect 418988 3256 419040 3262
rect 418988 3198 419040 3204
rect 416780 3188 416832 3194
rect 416780 3130 416832 3136
rect 417884 3052 417936 3058
rect 417884 2994 417936 3000
rect 417896 480 417924 2994
rect 419000 480 419028 3198
rect 420196 480 420224 4762
rect 420932 2990 420960 299338
rect 421024 6254 421052 301838
rect 421392 301838 421682 301866
rect 422312 301838 422510 301866
rect 421392 299402 421420 301838
rect 421380 299396 421432 299402
rect 421380 299338 421432 299344
rect 421012 6248 421064 6254
rect 421012 6190 421064 6196
rect 422312 4554 422340 301838
rect 423324 297430 423352 301852
rect 424152 298926 424180 301852
rect 424244 301838 424994 301866
rect 425072 301838 425822 301866
rect 426452 301838 426558 301866
rect 426636 301838 427386 301866
rect 427924 301838 428214 301866
rect 424140 298920 424192 298926
rect 424140 298862 424192 298868
rect 423588 298240 423640 298246
rect 423588 298182 423640 298188
rect 423312 297424 423364 297430
rect 423312 297366 423364 297372
rect 422300 4548 422352 4554
rect 422300 4490 422352 4496
rect 423600 3534 423628 298182
rect 424244 296714 424272 301838
rect 424968 298852 425020 298858
rect 424968 298794 425020 298800
rect 424324 298308 424376 298314
rect 424324 298250 424376 298256
rect 423784 296686 424272 296714
rect 423784 4486 423812 296686
rect 423772 4480 423824 4486
rect 423772 4422 423824 4428
rect 422576 3528 422628 3534
rect 422576 3470 422628 3476
rect 423588 3528 423640 3534
rect 423588 3470 423640 3476
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 421380 3460 421432 3466
rect 421380 3402 421432 3408
rect 420920 2984 420972 2990
rect 420920 2926 420972 2932
rect 421392 480 421420 3402
rect 422588 480 422616 3470
rect 423784 480 423812 3470
rect 424336 3466 424364 298250
rect 424324 3460 424376 3466
rect 424324 3402 424376 3408
rect 424980 480 425008 298794
rect 425072 11830 425100 301838
rect 425704 297424 425756 297430
rect 425704 297366 425756 297372
rect 425060 11824 425112 11830
rect 425060 11766 425112 11772
rect 425716 3534 425744 297366
rect 425704 3528 425756 3534
rect 425704 3470 425756 3476
rect 426164 3460 426216 3466
rect 426164 3402 426216 3408
rect 426176 480 426204 3402
rect 426452 3194 426480 301838
rect 426636 296714 426664 301838
rect 426544 296686 426664 296714
rect 426544 4418 426572 296686
rect 427924 11898 427952 301838
rect 429028 299266 429056 301852
rect 429212 301838 429870 301866
rect 430606 301838 430712 301866
rect 429016 299260 429068 299266
rect 429016 299202 429068 299208
rect 428464 297288 428516 297294
rect 428464 297230 428516 297236
rect 427912 11892 427964 11898
rect 427912 11834 427964 11840
rect 426532 4412 426584 4418
rect 426532 4354 426584 4360
rect 428476 3534 428504 297230
rect 429212 4350 429240 301838
rect 430580 299260 430632 299266
rect 430580 299202 430632 299208
rect 430488 298920 430540 298926
rect 430488 298862 430540 298868
rect 429200 4344 429252 4350
rect 429200 4286 429252 4292
rect 430500 3534 430528 298862
rect 430592 3602 430620 299202
rect 430684 10402 430712 301838
rect 431144 301838 431434 301866
rect 431972 301838 432262 301866
rect 432340 301838 433090 301866
rect 431144 299266 431172 301838
rect 431132 299260 431184 299266
rect 431132 299202 431184 299208
rect 430672 10396 430724 10402
rect 430672 10338 430724 10344
rect 431972 4282 432000 301838
rect 432340 296714 432368 301838
rect 433904 298790 433932 301852
rect 433892 298784 433944 298790
rect 433892 298726 433944 298732
rect 432604 297220 432656 297226
rect 432604 297162 432656 297168
rect 432064 296686 432368 296714
rect 432064 296206 432092 296686
rect 432052 296200 432104 296206
rect 432052 296142 432104 296148
rect 431960 4276 432012 4282
rect 431960 4218 432012 4224
rect 432052 3800 432104 3806
rect 432052 3742 432104 3748
rect 430580 3596 430632 3602
rect 430580 3538 430632 3544
rect 430856 3596 430908 3602
rect 430856 3538 430908 3544
rect 427268 3528 427320 3534
rect 427268 3470 427320 3476
rect 428464 3528 428516 3534
rect 428464 3470 428516 3476
rect 429660 3528 429712 3534
rect 429660 3470 429712 3476
rect 430488 3528 430540 3534
rect 430488 3470 430540 3476
rect 426440 3188 426492 3194
rect 426440 3130 426492 3136
rect 427280 480 427308 3470
rect 428464 3188 428516 3194
rect 428464 3130 428516 3136
rect 428476 480 428504 3130
rect 429672 480 429700 3470
rect 430868 480 430896 3538
rect 432064 480 432092 3742
rect 432616 3602 432644 297162
rect 434732 6662 434760 301852
rect 434824 301838 435482 301866
rect 434824 296138 434852 301838
rect 436296 299062 436324 301852
rect 436664 301838 437138 301866
rect 435364 299056 435416 299062
rect 435364 298998 435416 299004
rect 436284 299056 436336 299062
rect 436284 298998 436336 299004
rect 434812 296132 434864 296138
rect 434812 296074 434864 296080
rect 434720 6656 434772 6662
rect 434720 6598 434772 6604
rect 433248 3664 433300 3670
rect 433248 3606 433300 3612
rect 432604 3596 432656 3602
rect 432604 3538 432656 3544
rect 433260 480 433288 3606
rect 435376 3534 435404 298998
rect 436008 298240 436060 298246
rect 436008 298182 436060 298188
rect 436020 3534 436048 298182
rect 436664 296714 436692 301838
rect 437952 299062 437980 301852
rect 436744 299056 436796 299062
rect 436744 298998 436796 299004
rect 437940 299056 437992 299062
rect 437940 298998 437992 299004
rect 438124 299056 438176 299062
rect 438124 298998 438176 299004
rect 436204 296686 436692 296714
rect 436204 6730 436232 296686
rect 436756 7614 436784 298998
rect 436744 7608 436796 7614
rect 436744 7550 436796 7556
rect 436192 6724 436244 6730
rect 436192 6666 436244 6672
rect 437940 3596 437992 3602
rect 437940 3538 437992 3544
rect 435364 3528 435416 3534
rect 435364 3470 435416 3476
rect 435548 3528 435600 3534
rect 435548 3470 435600 3476
rect 436008 3528 436060 3534
rect 436008 3470 436060 3476
rect 436744 3528 436796 3534
rect 436744 3470 436796 3476
rect 434444 2848 434496 2854
rect 434444 2790 434496 2796
rect 434456 480 434484 2790
rect 435560 480 435588 3470
rect 436756 480 436784 3470
rect 437952 480 437980 3538
rect 438136 3534 438164 298998
rect 438780 298790 438808 301852
rect 438872 301838 439530 301866
rect 438768 298784 438820 298790
rect 438768 298726 438820 298732
rect 438872 6798 438900 301838
rect 440240 299532 440292 299538
rect 440240 299474 440292 299480
rect 439504 295996 439556 296002
rect 439504 295938 439556 295944
rect 438860 6792 438912 6798
rect 438860 6734 438912 6740
rect 439516 3602 439544 295938
rect 440252 3738 440280 299474
rect 440344 296070 440372 301852
rect 440896 301838 441186 301866
rect 440896 299538 440924 301838
rect 440884 299532 440936 299538
rect 440884 299474 440936 299480
rect 442000 297498 442028 301852
rect 442828 299130 442856 301852
rect 443288 301838 443670 301866
rect 442816 299124 442868 299130
rect 442816 299066 442868 299072
rect 442264 298988 442316 298994
rect 442264 298930 442316 298936
rect 441988 297492 442040 297498
rect 441988 297434 442040 297440
rect 440332 296064 440384 296070
rect 440332 296006 440384 296012
rect 441528 3800 441580 3806
rect 441528 3742 441580 3748
rect 440240 3732 440292 3738
rect 440240 3674 440292 3680
rect 440424 3664 440476 3670
rect 440424 3606 440476 3612
rect 439504 3596 439556 3602
rect 439504 3538 439556 3544
rect 438124 3528 438176 3534
rect 438124 3470 438176 3476
rect 439136 3052 439188 3058
rect 439136 2994 439188 3000
rect 439148 480 439176 2994
rect 440436 1850 440464 3606
rect 440344 1822 440464 1850
rect 440344 480 440372 1822
rect 441540 480 441568 3742
rect 442276 2990 442304 298930
rect 443288 298586 443316 301838
rect 443644 299124 443696 299130
rect 443644 299066 443696 299072
rect 443276 298580 443328 298586
rect 443276 298522 443328 298528
rect 443656 6390 443684 299066
rect 444288 298580 444340 298586
rect 444288 298522 444340 298528
rect 444300 6914 444328 298522
rect 444392 297566 444420 301852
rect 445220 299130 445248 301852
rect 445208 299124 445260 299130
rect 445208 299066 445260 299072
rect 446048 298994 446076 301852
rect 446140 301838 446890 301866
rect 446036 298988 446088 298994
rect 446036 298930 446088 298936
rect 444380 297560 444432 297566
rect 444380 297502 444432 297508
rect 446140 296714 446168 301838
rect 447704 298450 447732 301852
rect 447692 298444 447744 298450
rect 447692 298386 447744 298392
rect 447048 298240 447100 298246
rect 447048 298182 447100 298188
rect 443840 6886 444328 6914
rect 445864 296686 446168 296714
rect 443644 6384 443696 6390
rect 443644 6326 443696 6332
rect 442264 2984 442316 2990
rect 442264 2926 442316 2932
rect 442632 2984 442684 2990
rect 442632 2926 442684 2932
rect 442644 480 442672 2926
rect 443840 480 443868 6886
rect 445864 6322 445892 296686
rect 445852 6316 445904 6322
rect 445852 6258 445904 6264
rect 445024 3800 445076 3806
rect 445024 3742 445076 3748
rect 445036 480 445064 3742
rect 447060 3738 447088 298182
rect 448440 298178 448468 301852
rect 449164 299124 449216 299130
rect 449164 299066 449216 299072
rect 448428 298172 448480 298178
rect 448428 298114 448480 298120
rect 447784 297492 447836 297498
rect 447784 297434 447836 297440
rect 447796 3806 447824 297434
rect 447876 297152 447928 297158
rect 447876 297094 447928 297100
rect 447784 3800 447836 3806
rect 447784 3742 447836 3748
rect 446220 3732 446272 3738
rect 446220 3674 446272 3680
rect 447048 3732 447100 3738
rect 447048 3674 447100 3680
rect 447416 3732 447468 3738
rect 447416 3674 447468 3680
rect 446232 480 446260 3674
rect 447428 480 447456 3674
rect 447888 2854 447916 297094
rect 449176 6458 449204 299066
rect 449268 297634 449296 301852
rect 450096 299130 450124 301852
rect 450188 301838 450938 301866
rect 450084 299124 450136 299130
rect 450084 299066 450136 299072
rect 449808 298988 449860 298994
rect 449808 298930 449860 298936
rect 449256 297628 449308 297634
rect 449256 297570 449308 297576
rect 449164 6452 449216 6458
rect 449164 6394 449216 6400
rect 447876 2848 447928 2854
rect 447876 2790 447928 2796
rect 448612 2848 448664 2854
rect 448612 2790 448664 2796
rect 448624 480 448652 2790
rect 449820 480 449848 298930
rect 450188 296714 450216 301838
rect 451188 298580 451240 298586
rect 451188 298522 451240 298528
rect 450004 296686 450216 296714
rect 450004 3874 450032 296686
rect 451200 6914 451228 298522
rect 451752 297702 451780 301852
rect 452580 298518 452608 301852
rect 453316 298722 453344 301852
rect 453304 298716 453356 298722
rect 453304 298658 453356 298664
rect 452568 298512 452620 298518
rect 452568 298454 452620 298460
rect 454144 297770 454172 301852
rect 454236 301838 454986 301866
rect 455432 301838 455814 301866
rect 454132 297764 454184 297770
rect 454132 297706 454184 297712
rect 451740 297696 451792 297702
rect 451740 297638 451792 297644
rect 453304 297560 453356 297566
rect 453304 297502 453356 297508
rect 450924 6886 451228 6914
rect 449992 3868 450044 3874
rect 449992 3810 450044 3816
rect 450924 480 450952 6886
rect 453316 3330 453344 297502
rect 453396 297084 453448 297090
rect 453396 297026 453448 297032
rect 452108 3324 452160 3330
rect 452108 3266 452160 3272
rect 453304 3324 453356 3330
rect 453304 3266 453356 3272
rect 452120 480 452148 3266
rect 453408 3074 453436 297026
rect 454236 296714 454264 301838
rect 454052 296686 454264 296714
rect 454052 3942 454080 296686
rect 455432 4010 455460 301838
rect 456064 299192 456116 299198
rect 456064 299134 456116 299140
rect 455420 4004 455472 4010
rect 455420 3946 455472 3952
rect 454040 3936 454092 3942
rect 454040 3878 454092 3884
rect 454500 3936 454552 3942
rect 454500 3878 454552 3884
rect 453224 3046 453436 3074
rect 453224 2922 453252 3046
rect 453212 2916 453264 2922
rect 453212 2858 453264 2864
rect 453304 2916 453356 2922
rect 453304 2858 453356 2864
rect 453316 480 453344 2858
rect 454512 480 454540 3878
rect 456076 3738 456104 299134
rect 456628 297838 456656 301852
rect 457364 298722 457392 301852
rect 457352 298716 457404 298722
rect 457352 298658 457404 298664
rect 458192 298654 458220 301852
rect 458180 298648 458232 298654
rect 458180 298590 458232 298596
rect 458088 298512 458140 298518
rect 458088 298454 458140 298460
rect 456616 297832 456668 297838
rect 456616 297774 456668 297780
rect 457444 297628 457496 297634
rect 457444 297570 457496 297576
rect 456064 3732 456116 3738
rect 456064 3674 456116 3680
rect 456892 3732 456944 3738
rect 456892 3674 456944 3680
rect 455696 3324 455748 3330
rect 455696 3266 455748 3272
rect 455708 480 455736 3266
rect 456904 480 456932 3674
rect 457456 3330 457484 297570
rect 457444 3324 457496 3330
rect 457444 3266 457496 3272
rect 458100 480 458128 298454
rect 459020 297906 459048 301852
rect 459756 301838 459862 301866
rect 459008 297900 459060 297906
rect 459008 297842 459060 297848
rect 459192 4888 459244 4894
rect 459192 4830 459244 4836
rect 459204 480 459232 4830
rect 459756 4078 459784 301838
rect 460676 299198 460704 301852
rect 460664 299192 460716 299198
rect 460664 299134 460716 299140
rect 460204 298716 460256 298722
rect 460204 298658 460256 298664
rect 459744 4072 459796 4078
rect 459744 4014 459796 4020
rect 460216 3126 460244 298658
rect 461504 297974 461532 301852
rect 462240 298382 462268 301852
rect 463068 299334 463096 301852
rect 463056 299328 463108 299334
rect 463056 299270 463108 299276
rect 462228 298376 462280 298382
rect 462228 298318 462280 298324
rect 463896 298110 463924 301852
rect 463988 301838 464738 301866
rect 463884 298104 463936 298110
rect 463884 298046 463936 298052
rect 461492 297968 461544 297974
rect 461492 297910 461544 297916
rect 461584 297900 461636 297906
rect 461584 297842 461636 297848
rect 461596 6914 461624 297842
rect 463988 296714 464016 301838
rect 465552 298722 465580 301852
rect 465540 298716 465592 298722
rect 465540 298658 465592 298664
rect 465724 298512 465776 298518
rect 465724 298454 465776 298460
rect 464344 297696 464396 297702
rect 464344 297638 464396 297644
rect 461504 6886 461624 6914
rect 463712 296686 464016 296714
rect 460388 4004 460440 4010
rect 460388 3946 460440 3952
rect 460204 3120 460256 3126
rect 460204 3062 460256 3068
rect 460400 480 460428 3946
rect 461504 2854 461532 6886
rect 463712 4146 463740 296686
rect 463700 4140 463752 4146
rect 463700 4082 463752 4088
rect 461584 3868 461636 3874
rect 461584 3810 461636 3816
rect 461492 2848 461544 2854
rect 461492 2790 461544 2796
rect 461596 480 461624 3810
rect 464356 3398 464384 297638
rect 465736 3806 465764 298454
rect 466288 297362 466316 301852
rect 467116 299470 467144 301852
rect 467104 299464 467156 299470
rect 467104 299406 467156 299412
rect 467944 299402 467972 301852
rect 467932 299396 467984 299402
rect 467932 299338 467984 299344
rect 467748 299328 467800 299334
rect 467748 299270 467800 299276
rect 466368 298716 466420 298722
rect 466368 298658 466420 298664
rect 466276 297356 466328 297362
rect 466276 297298 466328 297304
rect 465724 3800 465776 3806
rect 465724 3742 465776 3748
rect 466380 3398 466408 298658
rect 467760 6914 467788 299270
rect 468772 298042 468800 301852
rect 469324 301838 469614 301866
rect 470152 301838 470442 301866
rect 470612 301838 471178 301866
rect 469220 299328 469272 299334
rect 469220 299270 469272 299276
rect 468760 298036 468812 298042
rect 468760 297978 468812 297984
rect 468484 297832 468536 297838
rect 468484 297774 468536 297780
rect 467484 6886 467788 6914
rect 462780 3392 462832 3398
rect 462780 3334 462832 3340
rect 464344 3392 464396 3398
rect 464344 3334 464396 3340
rect 465172 3392 465224 3398
rect 465172 3334 465224 3340
rect 466368 3392 466420 3398
rect 466368 3334 466420 3340
rect 462792 480 462820 3334
rect 463976 3120 464028 3126
rect 463976 3062 464028 3068
rect 463988 480 464016 3062
rect 465184 480 465212 3334
rect 466276 3324 466328 3330
rect 466276 3266 466328 3272
rect 466288 480 466316 3266
rect 467484 480 467512 6886
rect 468496 3330 468524 297774
rect 469232 4146 469260 299270
rect 469220 4140 469272 4146
rect 469220 4082 469272 4088
rect 468668 4072 468720 4078
rect 468668 4014 468720 4020
rect 468484 3324 468536 3330
rect 468484 3266 468536 3272
rect 468680 480 468708 4014
rect 469324 3262 469352 301838
rect 470152 299334 470180 301838
rect 470140 299328 470192 299334
rect 470140 299270 470192 299276
rect 470612 4826 470640 301838
rect 471992 298314 472020 301852
rect 472624 299396 472676 299402
rect 472624 299338 472676 299344
rect 471980 298308 472032 298314
rect 471980 298250 472032 298256
rect 471244 297764 471296 297770
rect 471244 297706 471296 297712
rect 470600 4820 470652 4826
rect 470600 4762 470652 4768
rect 471256 4146 471284 297706
rect 469864 4140 469916 4146
rect 469864 4082 469916 4088
rect 471244 4140 471296 4146
rect 471244 4082 471296 4088
rect 469312 3256 469364 3262
rect 469312 3198 469364 3204
rect 469876 480 469904 4082
rect 472256 3800 472308 3806
rect 472256 3742 472308 3748
rect 471060 3528 471112 3534
rect 471060 3470 471112 3476
rect 471072 480 471100 3470
rect 472268 480 472296 3742
rect 472636 3194 472664 299338
rect 472820 298858 472848 301852
rect 472808 298852 472860 298858
rect 472808 298794 472860 298800
rect 473648 297430 473676 301852
rect 474004 299464 474056 299470
rect 474004 299406 474056 299412
rect 473636 297424 473688 297430
rect 473636 297366 473688 297372
rect 474016 3602 474044 299406
rect 474476 298926 474504 301852
rect 474752 301838 475318 301866
rect 474464 298920 474516 298926
rect 474464 298862 474516 298868
rect 474096 298444 474148 298450
rect 474096 298386 474148 298392
rect 474004 3596 474056 3602
rect 474004 3538 474056 3544
rect 472624 3188 472676 3194
rect 472624 3130 472676 3136
rect 473452 3188 473504 3194
rect 473452 3130 473504 3136
rect 473464 480 473492 3130
rect 474108 3058 474136 298386
rect 474752 3466 474780 301838
rect 475384 298852 475436 298858
rect 475384 298794 475436 298800
rect 474740 3460 474792 3466
rect 474740 3402 474792 3408
rect 474556 3256 474608 3262
rect 474556 3198 474608 3204
rect 474096 3052 474148 3058
rect 474096 2994 474148 3000
rect 474568 480 474596 3198
rect 475396 2922 475424 298794
rect 476040 297294 476068 301852
rect 476868 299402 476896 301852
rect 476856 299396 476908 299402
rect 476856 299338 476908 299344
rect 477696 299266 477724 301852
rect 478144 299396 478196 299402
rect 478144 299338 478196 299344
rect 477684 299260 477736 299266
rect 477684 299202 477736 299208
rect 476764 298920 476816 298926
rect 476764 298862 476816 298868
rect 476028 297288 476080 297294
rect 476028 297230 476080 297236
rect 475752 4072 475804 4078
rect 475752 4014 475804 4020
rect 475384 2916 475436 2922
rect 475384 2858 475436 2864
rect 475764 480 475792 4014
rect 476776 2990 476804 298862
rect 478156 6914 478184 299338
rect 478236 299260 478288 299266
rect 478236 299202 478288 299208
rect 478064 6886 478184 6914
rect 478064 3534 478092 6886
rect 478052 3528 478104 3534
rect 478052 3470 478104 3476
rect 478248 3466 478276 299202
rect 478524 297226 478552 301852
rect 479352 299470 479380 301852
rect 479340 299464 479392 299470
rect 479340 299406 479392 299412
rect 480088 299266 480116 301852
rect 480640 301838 480930 301866
rect 480076 299260 480128 299266
rect 480076 299202 480128 299208
rect 480168 299260 480220 299266
rect 480168 299202 480220 299208
rect 480180 299010 480208 299202
rect 480088 298982 480208 299010
rect 480088 298178 480116 298982
rect 480168 298852 480220 298858
rect 480168 298794 480220 298800
rect 479524 298172 479576 298178
rect 479524 298114 479576 298120
rect 480076 298172 480128 298178
rect 480076 298114 480128 298120
rect 478512 297220 478564 297226
rect 478512 297162 478564 297168
rect 479536 3670 479564 298114
rect 479524 3664 479576 3670
rect 479524 3606 479576 3612
rect 480180 3534 480208 298794
rect 480640 297158 480668 301838
rect 481744 298790 481772 301852
rect 482572 299062 482600 301852
rect 483124 301838 483414 301866
rect 482560 299056 482612 299062
rect 482560 298998 482612 299004
rect 481732 298784 481784 298790
rect 481732 298726 481784 298732
rect 482928 298784 482980 298790
rect 482928 298726 482980 298732
rect 482284 298648 482336 298654
rect 482284 298590 482336 298596
rect 480904 298308 480956 298314
rect 480904 298250 480956 298256
rect 480628 297152 480680 297158
rect 480628 297094 480680 297100
rect 480916 3942 480944 298250
rect 480904 3936 480956 3942
rect 480904 3878 480956 3884
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 480168 3528 480220 3534
rect 480168 3470 480220 3476
rect 478236 3460 478288 3466
rect 478236 3402 478288 3408
rect 478144 3392 478196 3398
rect 478144 3334 478196 3340
rect 476948 3324 477000 3330
rect 476948 3266 477000 3272
rect 476764 2984 476816 2990
rect 476764 2926 476816 2932
rect 476960 480 476988 3266
rect 478156 480 478184 3334
rect 479352 480 479380 3470
rect 481732 3460 481784 3466
rect 481732 3402 481784 3408
rect 480536 3256 480588 3262
rect 480536 3198 480588 3204
rect 480548 480 480576 3198
rect 481744 480 481772 3402
rect 482296 3194 482324 298590
rect 482836 3528 482888 3534
rect 482836 3470 482888 3476
rect 482284 3188 482336 3194
rect 482284 3130 482336 3136
rect 482848 480 482876 3470
rect 482940 3466 482968 298726
rect 483124 296002 483152 301838
rect 484228 298450 484256 301852
rect 484964 299266 484992 301852
rect 484952 299260 485004 299266
rect 484952 299202 485004 299208
rect 485688 299056 485740 299062
rect 485688 298998 485740 299004
rect 484216 298444 484268 298450
rect 484216 298386 484268 298392
rect 483664 298376 483716 298382
rect 483664 298318 483716 298324
rect 483112 295996 483164 296002
rect 483112 295938 483164 295944
rect 482928 3460 482980 3466
rect 482928 3402 482980 3408
rect 483676 3126 483704 298318
rect 484308 297424 484360 297430
rect 484308 297366 484360 297372
rect 484320 6914 484348 297366
rect 484044 6886 484348 6914
rect 483664 3120 483716 3126
rect 483664 3062 483716 3068
rect 484044 480 484072 6886
rect 485700 3534 485728 298998
rect 485792 297090 485820 301852
rect 486620 298926 486648 301852
rect 487448 298994 487476 301852
rect 487436 298988 487488 298994
rect 487436 298930 487488 298936
rect 486608 298920 486660 298926
rect 486608 298862 486660 298868
rect 487068 298920 487120 298926
rect 487068 298862 487120 298868
rect 486424 298172 486476 298178
rect 486424 298114 486476 298120
rect 485780 297084 485832 297090
rect 485780 297026 485832 297032
rect 486436 6914 486464 298114
rect 486344 6886 486464 6914
rect 486344 4010 486372 6886
rect 486332 4004 486384 4010
rect 486332 3946 486384 3952
rect 485228 3528 485280 3534
rect 485228 3470 485280 3476
rect 485688 3528 485740 3534
rect 485688 3470 485740 3476
rect 485240 480 485268 3470
rect 487080 3058 487108 298862
rect 487804 298444 487856 298450
rect 487804 298386 487856 298392
rect 487816 3602 487844 298386
rect 488276 297498 488304 301852
rect 489012 298246 489040 301852
rect 489472 301838 489854 301866
rect 489472 298518 489500 301838
rect 489828 298988 489880 298994
rect 489828 298930 489880 298936
rect 489460 298512 489512 298518
rect 489460 298454 489512 298460
rect 489000 298240 489052 298246
rect 489000 298182 489052 298188
rect 489184 297968 489236 297974
rect 489184 297910 489236 297916
rect 488264 297492 488316 297498
rect 488264 297434 488316 297440
rect 487804 3596 487856 3602
rect 487804 3538 487856 3544
rect 488816 3596 488868 3602
rect 488816 3538 488868 3544
rect 487620 3528 487672 3534
rect 487620 3470 487672 3476
rect 486424 3052 486476 3058
rect 486424 2994 486476 3000
rect 487068 3052 487120 3058
rect 487068 2994 487120 3000
rect 486436 480 486464 2994
rect 487632 480 487660 3470
rect 488828 480 488856 3538
rect 489196 3534 489224 297910
rect 489840 3602 489868 298930
rect 490668 297906 490696 301852
rect 491496 299130 491524 301852
rect 491484 299124 491536 299130
rect 491484 299066 491536 299072
rect 492324 298586 492352 301852
rect 492312 298580 492364 298586
rect 492312 298522 492364 298528
rect 491944 298512 491996 298518
rect 491944 298454 491996 298460
rect 491208 298376 491260 298382
rect 491208 298318 491260 298324
rect 490656 297900 490708 297906
rect 490656 297842 490708 297848
rect 491116 297492 491168 297498
rect 491116 297434 491168 297440
rect 489828 3596 489880 3602
rect 489828 3538 489880 3544
rect 489920 3596 489972 3602
rect 489920 3538 489972 3544
rect 489184 3528 489236 3534
rect 489184 3470 489236 3476
rect 489932 480 489960 3538
rect 491128 480 491156 297434
rect 491220 3602 491248 298318
rect 491956 3874 491984 298454
rect 492036 298172 492088 298178
rect 492036 298114 492088 298120
rect 492048 3942 492076 298114
rect 493152 297566 493180 301852
rect 493888 299470 493916 301852
rect 493876 299464 493928 299470
rect 493876 299406 493928 299412
rect 493324 299260 493376 299266
rect 493324 299202 493376 299208
rect 493140 297560 493192 297566
rect 493140 297502 493192 297508
rect 492036 3936 492088 3942
rect 492036 3878 492088 3884
rect 491944 3868 491996 3874
rect 491944 3810 491996 3816
rect 493336 3738 493364 299202
rect 493968 299124 494020 299130
rect 493968 299066 494020 299072
rect 493324 3732 493376 3738
rect 493324 3674 493376 3680
rect 492312 3664 492364 3670
rect 492312 3606 492364 3612
rect 491208 3596 491260 3602
rect 491208 3538 491260 3544
rect 492324 480 492352 3606
rect 493980 3602 494008 299066
rect 494716 298314 494744 301852
rect 494704 298308 494756 298314
rect 494704 298250 494756 298256
rect 495544 297634 495572 301852
rect 496372 299266 496400 301852
rect 496360 299260 496412 299266
rect 496360 299202 496412 299208
rect 497200 299198 497228 301852
rect 497384 301838 497950 301866
rect 497188 299192 497240 299198
rect 497188 299134 497240 299140
rect 496728 298376 496780 298382
rect 496728 298318 496780 298324
rect 495532 297628 495584 297634
rect 495532 297570 495584 297576
rect 495348 297560 495400 297566
rect 495348 297502 495400 297508
rect 493508 3596 493560 3602
rect 493508 3538 493560 3544
rect 493968 3596 494020 3602
rect 493968 3538 494020 3544
rect 493520 480 493548 3538
rect 495360 3058 495388 297502
rect 496740 3602 496768 298318
rect 497384 296714 497412 301838
rect 497464 298512 497516 298518
rect 497464 298454 497516 298460
rect 496924 296686 497412 296714
rect 496924 4894 496952 296686
rect 496912 4888 496964 4894
rect 496912 4830 496964 4836
rect 497096 3868 497148 3874
rect 497096 3810 497148 3816
rect 495900 3596 495952 3602
rect 495900 3538 495952 3544
rect 496728 3596 496780 3602
rect 496728 3538 496780 3544
rect 494704 3052 494756 3058
rect 494704 2994 494756 3000
rect 495348 3052 495400 3058
rect 495348 2994 495400 3000
rect 494716 480 494744 2994
rect 495912 480 495940 3538
rect 497108 480 497136 3810
rect 497476 3330 497504 298454
rect 498764 298246 498792 301852
rect 499592 298586 499620 301852
rect 499580 298580 499632 298586
rect 499580 298522 499632 298528
rect 500224 298308 500276 298314
rect 500224 298250 500276 298256
rect 498752 298240 498804 298246
rect 498752 298182 498804 298188
rect 500236 4078 500264 298250
rect 500420 297702 500448 301852
rect 501248 299470 501276 301852
rect 501236 299464 501288 299470
rect 501236 299406 501288 299412
rect 502076 298722 502104 301852
rect 502064 298716 502116 298722
rect 502064 298658 502116 298664
rect 500868 298444 500920 298450
rect 500868 298386 500920 298392
rect 500408 297696 500460 297702
rect 500408 297638 500460 297644
rect 500880 6914 500908 298386
rect 501604 298376 501656 298382
rect 501604 298318 501656 298324
rect 500604 6886 500908 6914
rect 500224 4072 500276 4078
rect 500224 4014 500276 4020
rect 499396 3732 499448 3738
rect 499396 3674 499448 3680
rect 498200 3664 498252 3670
rect 498200 3606 498252 3612
rect 497464 3324 497516 3330
rect 497464 3266 497516 3272
rect 498212 480 498240 3606
rect 499408 480 499436 3674
rect 500604 480 500632 6886
rect 501616 3398 501644 298318
rect 502812 297838 502840 301852
rect 503640 299334 503668 301852
rect 503628 299328 503680 299334
rect 503628 299270 503680 299276
rect 504364 299328 504416 299334
rect 504364 299270 504416 299276
rect 503628 299192 503680 299198
rect 503628 299134 503680 299140
rect 502984 298580 503036 298586
rect 502984 298522 503036 298528
rect 502800 297832 502852 297838
rect 502800 297774 502852 297780
rect 501788 6180 501840 6186
rect 501788 6122 501840 6128
rect 501604 3392 501656 3398
rect 501604 3334 501656 3340
rect 501800 480 501828 6122
rect 502996 3738 503024 298522
rect 502984 3732 503036 3738
rect 502984 3674 503036 3680
rect 503640 3534 503668 299134
rect 504180 3936 504232 3942
rect 504180 3878 504232 3884
rect 502984 3528 503036 3534
rect 502984 3470 503036 3476
rect 503628 3528 503680 3534
rect 503628 3470 503680 3476
rect 502996 480 503024 3470
rect 504192 480 504220 3878
rect 504376 3806 504404 299270
rect 504468 298246 504496 301852
rect 504456 298240 504508 298246
rect 504456 298182 504508 298188
rect 505296 297770 505324 301852
rect 506124 299402 506152 301852
rect 506112 299396 506164 299402
rect 506112 299338 506164 299344
rect 506860 299334 506888 301852
rect 506848 299328 506900 299334
rect 506848 299270 506900 299276
rect 507688 298654 507716 301852
rect 508240 301838 508530 301866
rect 507768 299396 507820 299402
rect 507768 299338 507820 299344
rect 507676 298648 507728 298654
rect 507676 298590 507728 298596
rect 505284 297764 505336 297770
rect 505284 297706 505336 297712
rect 505376 4140 505428 4146
rect 505376 4082 505428 4088
rect 504364 3800 504416 3806
rect 504364 3742 504416 3748
rect 505388 480 505416 4082
rect 507676 3732 507728 3738
rect 507676 3674 507728 3680
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 506492 480 506520 3470
rect 507688 480 507716 3674
rect 507780 3534 507808 299338
rect 508240 298178 508268 301838
rect 509148 298716 509200 298722
rect 509148 298658 509200 298664
rect 508504 298444 508556 298450
rect 508504 298386 508556 298392
rect 508228 298172 508280 298178
rect 508228 298114 508280 298120
rect 507768 3528 507820 3534
rect 507768 3470 507820 3476
rect 508516 3398 508544 298386
rect 509160 6914 509188 298658
rect 509344 298314 509372 301852
rect 510172 298518 510200 301852
rect 510160 298512 510212 298518
rect 510160 298454 510212 298460
rect 511000 298382 511028 301852
rect 511736 298858 511764 301852
rect 512104 301838 512578 301866
rect 511724 298852 511776 298858
rect 511724 298794 511776 298800
rect 511908 298648 511960 298654
rect 511908 298590 511960 298596
rect 510988 298376 511040 298382
rect 510988 298318 511040 298324
rect 509332 298308 509384 298314
rect 509332 298250 509384 298256
rect 511264 298308 511316 298314
rect 511264 298250 511316 298256
rect 511276 6914 511304 298250
rect 508884 6886 509188 6914
rect 511184 6886 511304 6914
rect 508504 3392 508556 3398
rect 508504 3334 508556 3340
rect 508884 480 508912 6886
rect 511184 4146 511212 6886
rect 511172 4140 511224 4146
rect 511172 4082 511224 4088
rect 510068 3596 510120 3602
rect 510068 3538 510120 3544
rect 510080 480 510108 3538
rect 511920 3534 511948 298590
rect 511264 3528 511316 3534
rect 511264 3470 511316 3476
rect 511908 3528 511960 3534
rect 511908 3470 511960 3476
rect 511276 480 511304 3470
rect 512104 3466 512132 301838
rect 513288 298852 513340 298858
rect 513288 298794 513340 298800
rect 513300 3534 513328 298794
rect 513392 298790 513420 301852
rect 513380 298784 513432 298790
rect 513380 298726 513432 298732
rect 514220 298450 514248 301852
rect 514208 298444 514260 298450
rect 514208 298386 514260 298392
rect 515048 297430 515076 301852
rect 515324 301838 515798 301866
rect 515324 299062 515352 301838
rect 515312 299056 515364 299062
rect 515312 298998 515364 299004
rect 515404 299056 515456 299062
rect 515404 298998 515456 299004
rect 515036 297424 515088 297430
rect 515036 297366 515088 297372
rect 515416 3534 515444 298998
rect 516612 298926 516640 301852
rect 517072 301838 517454 301866
rect 516600 298920 516652 298926
rect 516600 298862 516652 298868
rect 516048 298784 516100 298790
rect 516048 298726 516100 298732
rect 516060 6914 516088 298726
rect 517072 297974 517100 301838
rect 518268 298994 518296 301852
rect 519096 299266 519124 301852
rect 519084 299260 519136 299266
rect 519084 299202 519136 299208
rect 519544 299260 519596 299266
rect 519544 299202 519596 299208
rect 518256 298988 518308 298994
rect 518256 298930 518308 298936
rect 518808 298988 518860 298994
rect 518808 298930 518860 298936
rect 517428 298920 517480 298926
rect 517428 298862 517480 298868
rect 517060 297968 517112 297974
rect 517060 297910 517112 297916
rect 517440 6914 517468 298862
rect 518164 298172 518216 298178
rect 518164 298114 518216 298120
rect 515968 6886 516088 6914
rect 517164 6886 517468 6914
rect 512460 3528 512512 3534
rect 512460 3470 512512 3476
rect 513288 3528 513340 3534
rect 513288 3470 513340 3476
rect 513564 3528 513616 3534
rect 513564 3470 513616 3476
rect 515404 3528 515456 3534
rect 515404 3470 515456 3476
rect 512092 3460 512144 3466
rect 512092 3402 512144 3408
rect 512472 480 512500 3470
rect 513576 480 513604 3470
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 514772 480 514800 3402
rect 515968 480 515996 6886
rect 517164 480 517192 6886
rect 518176 3806 518204 298114
rect 518164 3800 518216 3806
rect 518164 3742 518216 3748
rect 518820 3534 518848 298930
rect 519556 6914 519584 299202
rect 519924 297498 519952 301852
rect 520188 298444 520240 298450
rect 520188 298386 520240 298392
rect 519912 297492 519964 297498
rect 519912 297434 519964 297440
rect 519464 6886 519584 6914
rect 519464 3874 519492 6886
rect 519452 3868 519504 3874
rect 519452 3810 519504 3816
rect 520200 3534 520228 298386
rect 520660 298178 520688 301852
rect 521488 299130 521516 301852
rect 522040 301838 522330 301866
rect 521476 299124 521528 299130
rect 521476 299066 521528 299072
rect 521568 298580 521620 298586
rect 521568 298522 521620 298528
rect 520648 298172 520700 298178
rect 520648 298114 520700 298120
rect 521580 3534 521608 298522
rect 522040 297566 522068 301838
rect 523144 299470 523172 301852
rect 523132 299464 523184 299470
rect 523132 299406 523184 299412
rect 522396 299328 522448 299334
rect 522396 299270 522448 299276
rect 522304 298240 522356 298246
rect 522304 298182 522356 298188
rect 522028 297560 522080 297566
rect 522028 297502 522080 297508
rect 522316 3942 522344 298182
rect 522304 3936 522356 3942
rect 522304 3878 522356 3884
rect 521844 3800 521896 3806
rect 521844 3742 521896 3748
rect 518348 3528 518400 3534
rect 518348 3470 518400 3476
rect 518808 3528 518860 3534
rect 518808 3470 518860 3476
rect 519544 3528 519596 3534
rect 519544 3470 519596 3476
rect 520188 3528 520240 3534
rect 520188 3470 520240 3476
rect 520740 3528 520792 3534
rect 520740 3470 520792 3476
rect 521568 3528 521620 3534
rect 521568 3470 521620 3476
rect 518360 480 518388 3470
rect 519556 480 519584 3470
rect 520752 480 520780 3470
rect 521856 480 521884 3742
rect 522408 3670 522436 299270
rect 523972 299266 524000 301852
rect 524708 299334 524736 301852
rect 524696 299328 524748 299334
rect 524696 299270 524748 299276
rect 525156 299328 525208 299334
rect 525156 299270 525208 299276
rect 523960 299260 524012 299266
rect 523960 299202 524012 299208
rect 525064 298444 525116 298450
rect 525064 298386 525116 298392
rect 524236 4072 524288 4078
rect 524236 4014 524288 4020
rect 522396 3664 522448 3670
rect 522396 3606 522448 3612
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523052 480 523080 3470
rect 524248 480 524276 4014
rect 525076 3602 525104 298386
rect 525168 6186 525196 299270
rect 525536 298518 525564 301852
rect 526364 299198 526392 301852
rect 526444 299464 526496 299470
rect 526444 299406 526496 299412
rect 526352 299192 526404 299198
rect 526352 299134 526404 299140
rect 525524 298512 525576 298518
rect 525524 298454 525576 298460
rect 525156 6180 525208 6186
rect 525156 6122 525208 6128
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 525432 3596 525484 3602
rect 525432 3538 525484 3544
rect 525444 480 525472 3538
rect 526456 3534 526484 299406
rect 527192 299334 527220 301852
rect 527180 299328 527232 299334
rect 527180 299270 527232 299276
rect 527088 299192 527140 299198
rect 527088 299134 527140 299140
rect 527100 3534 527128 299134
rect 528020 299130 528048 301852
rect 528008 299124 528060 299130
rect 528008 299066 528060 299072
rect 528848 298246 528876 301852
rect 529296 299328 529348 299334
rect 529296 299270 529348 299276
rect 529204 298580 529256 298586
rect 529204 298522 529256 298528
rect 528836 298240 528888 298246
rect 528836 298182 528888 298188
rect 529216 4078 529244 298522
rect 529204 4072 529256 4078
rect 529204 4014 529256 4020
rect 529308 3738 529336 299270
rect 529584 298314 529612 301852
rect 530412 299402 530440 301852
rect 530400 299396 530452 299402
rect 530400 299338 530452 299344
rect 530584 299396 530636 299402
rect 530584 299338 530636 299344
rect 529572 298308 529624 298314
rect 529572 298250 529624 298256
rect 529296 3732 529348 3738
rect 529296 3674 529348 3680
rect 526444 3528 526496 3534
rect 526444 3470 526496 3476
rect 526628 3528 526680 3534
rect 526628 3470 526680 3476
rect 527088 3528 527140 3534
rect 527088 3470 527140 3476
rect 527824 3528 527876 3534
rect 527824 3470 527876 3476
rect 526640 480 526668 3470
rect 527836 480 527864 3470
rect 530596 3466 530624 299338
rect 531240 299334 531268 301852
rect 531228 299328 531280 299334
rect 531228 299270 531280 299276
rect 531228 298920 531280 298926
rect 531228 298862 531280 298868
rect 530584 3460 530636 3466
rect 530584 3402 530636 3408
rect 531240 3398 531268 298862
rect 532068 298722 532096 301852
rect 532056 298716 532108 298722
rect 532056 298658 532108 298664
rect 532896 298450 532924 301852
rect 533724 298722 533752 301852
rect 533988 299328 534040 299334
rect 533988 299270 534040 299276
rect 533712 298716 533764 298722
rect 533712 298658 533764 298664
rect 533344 298648 533396 298654
rect 533344 298590 533396 298596
rect 532884 298444 532936 298450
rect 532884 298386 532936 298392
rect 531320 3868 531372 3874
rect 531320 3810 531372 3816
rect 530124 3392 530176 3398
rect 530124 3334 530176 3340
rect 531228 3392 531280 3398
rect 531228 3334 531280 3340
rect 529020 3324 529072 3330
rect 529020 3266 529072 3272
rect 529032 480 529060 3266
rect 530136 480 530164 3334
rect 531332 480 531360 3810
rect 533356 3806 533384 298590
rect 534000 6914 534028 299270
rect 534460 298858 534488 301852
rect 535288 299062 535316 301852
rect 536116 299402 536144 301852
rect 536104 299396 536156 299402
rect 536104 299338 536156 299344
rect 535276 299056 535328 299062
rect 535276 298998 535328 299004
rect 536196 299056 536248 299062
rect 536196 298998 536248 299004
rect 534448 298852 534500 298858
rect 534448 298794 534500 298800
rect 535368 298852 535420 298858
rect 535368 298794 535420 298800
rect 533724 6886 534028 6914
rect 533344 3800 533396 3806
rect 533344 3742 533396 3748
rect 532516 3188 532568 3194
rect 532516 3130 532568 3136
rect 532528 480 532556 3130
rect 533724 480 533752 6886
rect 535380 3534 535408 298794
rect 536104 298444 536156 298450
rect 536104 298386 536156 298392
rect 536116 3602 536144 298386
rect 536208 3738 536236 298998
rect 536944 298518 536972 301852
rect 537772 298790 537800 301852
rect 538508 298994 538536 301852
rect 539336 299266 539364 301852
rect 539324 299260 539376 299266
rect 539324 299202 539376 299208
rect 540164 299130 540192 301852
rect 540244 299260 540296 299266
rect 540244 299202 540296 299208
rect 540152 299124 540204 299130
rect 540152 299066 540204 299072
rect 538496 298988 538548 298994
rect 538496 298930 538548 298936
rect 538128 298920 538180 298926
rect 538128 298862 538180 298868
rect 537760 298784 537812 298790
rect 537760 298726 537812 298732
rect 536932 298512 536984 298518
rect 536932 298454 536984 298460
rect 537484 298512 537536 298518
rect 537484 298454 537536 298460
rect 536196 3732 536248 3738
rect 536196 3674 536248 3680
rect 536104 3596 536156 3602
rect 536104 3538 536156 3544
rect 534908 3528 534960 3534
rect 534908 3470 534960 3476
rect 535368 3528 535420 3534
rect 535368 3470 535420 3476
rect 537208 3528 537260 3534
rect 537208 3470 537260 3476
rect 534920 480 534948 3470
rect 536104 3392 536156 3398
rect 536104 3334 536156 3340
rect 536116 480 536144 3334
rect 537220 480 537248 3470
rect 537496 3330 537524 298454
rect 538140 3534 538168 298862
rect 539508 298784 539560 298790
rect 539508 298726 539560 298732
rect 538864 298716 538916 298722
rect 538864 298658 538916 298664
rect 538128 3528 538180 3534
rect 538128 3470 538180 3476
rect 538404 3528 538456 3534
rect 538404 3470 538456 3476
rect 537484 3324 537536 3330
rect 537484 3266 537536 3272
rect 538416 480 538444 3470
rect 538876 3194 538904 298658
rect 539520 3534 539548 298726
rect 539508 3528 539560 3534
rect 539508 3470 539560 3476
rect 540256 3398 540284 299202
rect 540888 298988 540940 298994
rect 540888 298930 540940 298936
rect 540900 6914 540928 298930
rect 540992 298654 541020 301852
rect 541820 299470 541848 301852
rect 541808 299464 541860 299470
rect 541808 299406 541860 299412
rect 540980 298648 541032 298654
rect 540980 298590 541032 298596
rect 542648 298586 542676 301852
rect 543384 299130 543412 301852
rect 544212 299198 544240 301852
rect 544672 301838 545054 301866
rect 544200 299192 544252 299198
rect 544200 299134 544252 299140
rect 544384 299192 544436 299198
rect 544384 299134 544436 299140
rect 543372 299124 543424 299130
rect 543372 299066 543424 299072
rect 543004 299056 543056 299062
rect 543004 298998 543056 299004
rect 542636 298580 542688 298586
rect 542636 298522 542688 298528
rect 540808 6886 540928 6914
rect 540244 3392 540296 3398
rect 540244 3334 540296 3340
rect 538864 3188 538916 3194
rect 538864 3130 538916 3136
rect 539600 3188 539652 3194
rect 539600 3130 539652 3136
rect 539612 480 539640 3130
rect 540808 480 540836 6886
rect 543016 3534 543044 298998
rect 543096 298648 543148 298654
rect 543096 298590 543148 298596
rect 541992 3528 542044 3534
rect 541992 3470 542044 3476
rect 543004 3528 543056 3534
rect 543004 3470 543056 3476
rect 542004 480 542032 3470
rect 543108 3194 543136 298590
rect 544396 3670 544424 299134
rect 544672 298450 544700 301838
rect 545028 299124 545080 299130
rect 545028 299066 545080 299072
rect 544660 298444 544712 298450
rect 544660 298386 544712 298392
rect 543188 3664 543240 3670
rect 543188 3606 543240 3612
rect 544384 3664 544436 3670
rect 544384 3606 544436 3612
rect 543096 3188 543148 3194
rect 543096 3130 543148 3136
rect 543200 480 543228 3606
rect 545040 3534 545068 299066
rect 545868 298518 545896 301852
rect 546696 299334 546724 301852
rect 546880 301838 547446 301866
rect 546684 299328 546736 299334
rect 546684 299270 546736 299276
rect 545856 298512 545908 298518
rect 545856 298454 545908 298460
rect 546880 296714 546908 301838
rect 547144 299464 547196 299470
rect 547144 299406 547196 299412
rect 546696 296686 546908 296714
rect 546696 3874 546724 296686
rect 546684 3868 546736 3874
rect 546684 3810 546736 3816
rect 546684 3732 546736 3738
rect 546684 3674 546736 3680
rect 544384 3528 544436 3534
rect 544384 3470 544436 3476
rect 545028 3528 545080 3534
rect 545028 3470 545080 3476
rect 545488 3528 545540 3534
rect 545488 3470 545540 3476
rect 544396 480 544424 3470
rect 545500 480 545528 3470
rect 546696 480 546724 3674
rect 547156 3534 547184 299406
rect 548260 298722 548288 301852
rect 549088 299402 549116 301852
rect 549076 299396 549128 299402
rect 549076 299338 549128 299344
rect 548524 299328 548576 299334
rect 548524 299270 548576 299276
rect 548248 298716 548300 298722
rect 548248 298658 548300 298664
rect 548536 3738 548564 299270
rect 549916 298858 549944 301852
rect 550744 299266 550772 301852
rect 550732 299260 550784 299266
rect 550732 299202 550784 299208
rect 551572 298926 551600 301852
rect 551928 299260 551980 299266
rect 551928 299202 551980 299208
rect 551560 298920 551612 298926
rect 551560 298862 551612 298868
rect 549904 298852 549956 298858
rect 549904 298794 549956 298800
rect 551284 298852 551336 298858
rect 551284 298794 551336 298800
rect 549168 298716 549220 298722
rect 549168 298658 549220 298664
rect 548524 3732 548576 3738
rect 548524 3674 548576 3680
rect 549076 3596 549128 3602
rect 549076 3538 549128 3544
rect 547144 3528 547196 3534
rect 547144 3470 547196 3476
rect 547880 3528 547932 3534
rect 547880 3470 547932 3476
rect 547892 480 547920 3470
rect 549088 480 549116 3538
rect 549180 3534 549208 298658
rect 551296 3534 551324 298794
rect 551940 3534 551968 299202
rect 552308 298790 552336 301852
rect 552296 298784 552348 298790
rect 552296 298726 552348 298732
rect 553136 298654 553164 301852
rect 553964 298994 553992 301852
rect 554792 299062 554820 301852
rect 555344 301838 555634 301866
rect 555344 299198 555372 301838
rect 555332 299192 555384 299198
rect 555332 299134 555384 299140
rect 555424 299192 555476 299198
rect 555424 299134 555476 299140
rect 554780 299056 554832 299062
rect 554780 298998 554832 299004
rect 553952 298988 554004 298994
rect 553952 298930 554004 298936
rect 553124 298648 553176 298654
rect 553124 298590 553176 298596
rect 554044 298172 554096 298178
rect 554044 298114 554096 298120
rect 554056 3602 554084 298114
rect 554044 3596 554096 3602
rect 554044 3538 554096 3544
rect 549168 3528 549220 3534
rect 549168 3470 549220 3476
rect 550272 3528 550324 3534
rect 550272 3470 550324 3476
rect 551284 3528 551336 3534
rect 551284 3470 551336 3476
rect 551468 3528 551520 3534
rect 551468 3470 551520 3476
rect 551928 3528 551980 3534
rect 551928 3470 551980 3476
rect 550284 480 550312 3470
rect 551480 480 551508 3470
rect 554964 3460 555016 3466
rect 554964 3402 555016 3408
rect 553768 3392 553820 3398
rect 553768 3334 553820 3340
rect 552664 3188 552716 3194
rect 552664 3130 552716 3136
rect 552676 480 552704 3130
rect 553780 480 553808 3334
rect 554976 480 555004 3402
rect 555436 3194 555464 299134
rect 556356 299130 556384 301852
rect 557184 299470 557212 301852
rect 557172 299464 557224 299470
rect 557172 299406 557224 299412
rect 558012 299334 558040 301852
rect 558184 299396 558236 299402
rect 558184 299338 558236 299344
rect 558000 299328 558052 299334
rect 558000 299270 558052 299276
rect 556344 299124 556396 299130
rect 556344 299066 556396 299072
rect 556804 298988 556856 298994
rect 556804 298930 556856 298936
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 555424 3188 555476 3194
rect 555424 3130 555476 3136
rect 556172 480 556200 3470
rect 556816 3466 556844 298930
rect 557448 298920 557500 298926
rect 557448 298862 557500 298868
rect 557460 3534 557488 298862
rect 557448 3528 557500 3534
rect 557448 3470 557500 3476
rect 556804 3460 556856 3466
rect 556804 3402 556856 3408
rect 558196 2990 558224 299338
rect 558840 298722 558868 301852
rect 558828 298716 558880 298722
rect 558828 298658 558880 298664
rect 558828 298580 558880 298586
rect 558828 298522 558880 298528
rect 558840 6914 558868 298522
rect 559668 298178 559696 301852
rect 560496 298858 560524 301852
rect 560944 299328 560996 299334
rect 560944 299270 560996 299276
rect 560484 298852 560536 298858
rect 560484 298794 560536 298800
rect 559656 298172 559708 298178
rect 559656 298114 559708 298120
rect 558564 6886 558868 6914
rect 557356 2984 557408 2990
rect 557356 2926 557408 2932
rect 558184 2984 558236 2990
rect 558184 2926 558236 2932
rect 557368 480 557396 2926
rect 558564 480 558592 6886
rect 560852 3528 560904 3534
rect 560852 3470 560904 3476
rect 559748 3460 559800 3466
rect 559748 3402 559800 3408
rect 559760 480 559788 3402
rect 560864 480 560892 3470
rect 560956 3466 560984 299270
rect 561232 299266 561260 301852
rect 561220 299260 561272 299266
rect 561220 299202 561272 299208
rect 562060 299198 562088 301852
rect 562244 301838 562902 301866
rect 562048 299192 562100 299198
rect 562048 299134 562100 299140
rect 561588 298308 561640 298314
rect 561588 298250 561640 298256
rect 561600 3534 561628 298250
rect 562244 296714 562272 301838
rect 563716 298994 563744 301852
rect 563704 298988 563756 298994
rect 563704 298930 563756 298936
rect 564544 298926 564572 301852
rect 565280 299402 565308 301852
rect 565268 299396 565320 299402
rect 565268 299338 565320 299344
rect 564532 298920 564584 298926
rect 564532 298862 564584 298868
rect 565728 298920 565780 298926
rect 565728 298862 565780 298868
rect 565084 298240 565136 298246
rect 565084 298182 565136 298188
rect 561876 296686 562272 296714
rect 561588 3528 561640 3534
rect 561588 3470 561640 3476
rect 560944 3460 560996 3466
rect 560944 3402 560996 3408
rect 561876 3398 561904 296686
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 561864 3392 561916 3398
rect 561864 3334 561916 3340
rect 562048 3324 562100 3330
rect 562048 3266 562100 3272
rect 562060 480 562088 3266
rect 563244 3188 563296 3194
rect 563244 3130 563296 3136
rect 563256 480 563284 3130
rect 564452 480 564480 3470
rect 565096 3194 565124 298182
rect 565636 3596 565688 3602
rect 565636 3538 565688 3544
rect 565084 3188 565136 3194
rect 565084 3130 565136 3136
rect 565648 480 565676 3538
rect 565740 3534 565768 298862
rect 566108 298586 566136 301852
rect 566936 299334 566964 301852
rect 566924 299328 566976 299334
rect 566924 299270 566976 299276
rect 567108 298784 567160 298790
rect 567108 298726 567160 298732
rect 566096 298580 566148 298586
rect 566096 298522 566148 298528
rect 566464 298172 566516 298178
rect 566464 298114 566516 298120
rect 565728 3528 565780 3534
rect 565728 3470 565780 3476
rect 566476 3330 566504 298114
rect 567120 6914 567148 298726
rect 567764 298314 567792 301852
rect 567752 298308 567804 298314
rect 567752 298250 567804 298256
rect 568592 298178 568620 301852
rect 569224 299396 569276 299402
rect 569224 299338 569276 299344
rect 568580 298172 568632 298178
rect 568580 298114 568632 298120
rect 566844 6886 567148 6914
rect 566464 3324 566516 3330
rect 566464 3266 566516 3272
rect 566844 480 566872 6886
rect 569236 3534 569264 299338
rect 569316 298716 569368 298722
rect 569316 298658 569368 298664
rect 569328 3602 569356 298658
rect 569420 298246 569448 301852
rect 570156 298926 570184 301852
rect 570144 298920 570196 298926
rect 570144 298862 570196 298868
rect 570984 298722 571012 301852
rect 571812 298790 571840 301852
rect 572640 299402 572668 301852
rect 572916 301838 573482 301866
rect 572628 299396 572680 299402
rect 572628 299338 572680 299344
rect 572628 299260 572680 299266
rect 572628 299202 572680 299208
rect 571800 298784 571852 298790
rect 571800 298726 571852 298732
rect 570972 298716 571024 298722
rect 570972 298658 571024 298664
rect 569408 298240 569460 298246
rect 569408 298182 569460 298188
rect 569316 3596 569368 3602
rect 569316 3538 569368 3544
rect 572640 3534 572668 299202
rect 568028 3528 568080 3534
rect 568028 3470 568080 3476
rect 569224 3528 569276 3534
rect 569224 3470 569276 3476
rect 571524 3528 571576 3534
rect 571524 3470 571576 3476
rect 572628 3528 572680 3534
rect 572628 3470 572680 3476
rect 568040 480 568068 3470
rect 570328 3460 570380 3466
rect 570328 3402 570380 3408
rect 569132 3256 569184 3262
rect 569132 3198 569184 3204
rect 569144 480 569172 3198
rect 570340 480 570368 3402
rect 571536 480 571564 3470
rect 572916 3262 572944 301838
rect 574008 299328 574060 299334
rect 574008 299270 574060 299276
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 572904 3256 572956 3262
rect 572904 3198 572956 3204
rect 572720 2916 572772 2922
rect 572720 2858 572772 2864
rect 572732 480 572760 2858
rect 573928 480 573956 3470
rect 574020 2922 574048 299270
rect 574204 3466 574232 301852
rect 575032 299266 575060 301852
rect 575860 299334 575888 301852
rect 576136 301838 576702 301866
rect 575848 299328 575900 299334
rect 575848 299270 575900 299276
rect 575020 299260 575072 299266
rect 575020 299202 575072 299208
rect 575388 298240 575440 298246
rect 575388 298182 575440 298188
rect 575400 6914 575428 298182
rect 576136 296714 576164 301838
rect 577516 298246 577544 301852
rect 577504 298240 577556 298246
rect 577504 298182 577556 298188
rect 578344 298178 578372 301852
rect 578436 301838 579094 301866
rect 579632 301838 579922 301866
rect 576768 298172 576820 298178
rect 576768 298114 576820 298120
rect 578332 298172 578384 298178
rect 578332 298114 578384 298120
rect 575124 6886 575428 6914
rect 575584 296686 576164 296714
rect 574192 3460 574244 3466
rect 574192 3402 574244 3408
rect 574008 2916 574060 2922
rect 574008 2858 574060 2864
rect 575124 480 575152 6886
rect 575584 3534 575612 296686
rect 576780 3534 576808 298114
rect 578436 3534 578464 301838
rect 575572 3528 575624 3534
rect 575572 3470 575624 3476
rect 576308 3528 576360 3534
rect 576308 3470 576360 3476
rect 576768 3528 576820 3534
rect 576768 3470 576820 3476
rect 577412 3528 577464 3534
rect 577412 3470 577464 3476
rect 578424 3528 578476 3534
rect 578424 3470 578476 3476
rect 576320 480 576348 3470
rect 577424 480 577452 3470
rect 579632 3058 579660 301838
rect 579804 139392 579856 139398
rect 579802 139360 579804 139369
rect 579856 139360 579858 139369
rect 579802 139295 579858 139304
rect 579988 113144 580040 113150
rect 579988 113086 580040 113092
rect 580000 112849 580028 113086
rect 579986 112840 580042 112849
rect 579986 112775 580042 112784
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 579802 33144 579858 33153
rect 579802 33079 579804 33088
rect 579856 33079 579858 33088
rect 579804 33050 579856 33056
rect 580172 20596 580224 20602
rect 580172 20538 580224 20544
rect 580184 19825 580212 20538
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 580276 6633 580304 302398
rect 580356 302388 580408 302394
rect 580356 302330 580408 302336
rect 580368 59673 580396 302330
rect 580750 301838 580856 301866
rect 580446 300112 580502 300121
rect 580446 300047 580502 300056
rect 580460 219065 580488 300047
rect 580446 219056 580502 219065
rect 580446 218991 580502 219000
rect 580354 59664 580410 59673
rect 580354 59599 580410 59608
rect 580828 16574 580856 301838
rect 581104 301838 581578 301866
rect 581104 16574 581132 301838
rect 582392 299334 582420 301852
rect 582380 299328 582432 299334
rect 582380 299270 582432 299276
rect 582484 232393 582512 702063
rect 583760 702024 583812 702030
rect 583760 701966 583812 701972
rect 583576 701888 583628 701894
rect 583576 701830 583628 701836
rect 582564 701820 582616 701826
rect 582564 701762 582616 701768
rect 582576 537849 582604 701762
rect 583392 701752 583444 701758
rect 583392 701694 583444 701700
rect 583208 701616 583260 701622
rect 583208 701558 583260 701564
rect 583116 701480 583168 701486
rect 583116 701422 583168 701428
rect 582932 701412 582984 701418
rect 582932 701354 582984 701360
rect 582748 700460 582800 700466
rect 582748 700402 582800 700408
rect 582654 700088 582710 700097
rect 582654 700023 582710 700032
rect 582562 537840 582618 537849
rect 582562 537775 582618 537784
rect 582668 272241 582696 700023
rect 582760 312089 582788 700402
rect 582840 700392 582892 700398
rect 582840 700334 582892 700340
rect 582852 325281 582880 700334
rect 582944 365129 582972 701354
rect 583024 701344 583076 701350
rect 583024 701286 583076 701292
rect 583036 378457 583064 701286
rect 583128 404977 583156 701422
rect 583220 418305 583248 701558
rect 583300 701548 583352 701554
rect 583300 701490 583352 701496
rect 583312 431633 583340 701490
rect 583404 471481 583432 701694
rect 583484 701684 583536 701690
rect 583484 701626 583536 701632
rect 583496 485217 583524 701626
rect 583588 525065 583616 701830
rect 583668 700528 583720 700534
rect 583668 700470 583720 700476
rect 583680 578241 583708 700470
rect 583772 631417 583800 701966
rect 583852 701956 583904 701962
rect 583852 701898 583904 701904
rect 583864 644337 583892 701898
rect 583850 644328 583906 644337
rect 583850 644263 583906 644272
rect 583758 631408 583814 631417
rect 583758 631343 583814 631352
rect 583758 579592 583814 579601
rect 583758 579527 583814 579536
rect 583666 578232 583722 578241
rect 583666 578167 583722 578176
rect 583574 525056 583630 525065
rect 583574 524991 583630 525000
rect 583482 485208 583538 485217
rect 583482 485143 583538 485152
rect 583390 471472 583446 471481
rect 583390 471407 583446 471416
rect 583298 431624 583354 431633
rect 583298 431559 583354 431568
rect 583206 418296 583262 418305
rect 583206 418231 583262 418240
rect 583114 404968 583170 404977
rect 583114 404903 583170 404912
rect 583022 378448 583078 378457
rect 583022 378383 583078 378392
rect 582930 365120 582986 365129
rect 582930 365055 582986 365064
rect 582838 325272 582894 325281
rect 582838 325207 582894 325216
rect 582746 312080 582802 312089
rect 582746 312015 582802 312024
rect 582748 298784 582800 298790
rect 582746 298752 582748 298761
rect 582800 298752 582802 298761
rect 582746 298687 582802 298696
rect 582654 272232 582710 272241
rect 582654 272167 582710 272176
rect 582656 258936 582708 258942
rect 582654 258904 582656 258913
rect 582708 258904 582710 258913
rect 582654 258839 582710 258848
rect 582470 232384 582526 232393
rect 582470 232319 582526 232328
rect 582564 165912 582616 165918
rect 582562 165880 582564 165889
rect 582616 165880 582618 165889
rect 582562 165815 582618 165824
rect 582472 152720 582524 152726
rect 582470 152688 582472 152697
rect 582524 152688 582526 152697
rect 582470 152623 582526 152632
rect 583772 20670 583800 579527
rect 583760 20664 583812 20670
rect 583760 20606 583812 20612
rect 580828 16546 580948 16574
rect 581104 16546 581776 16574
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 580920 3482 580948 16546
rect 580920 3454 581040 3482
rect 578608 3052 578660 3058
rect 578608 2994 578660 3000
rect 579620 3052 579672 3058
rect 579620 2994 579672 3000
rect 578620 480 578648 2994
rect 581012 480 581040 3454
rect 581748 490 581776 16546
rect 583392 3188 583444 3194
rect 583392 3130 583444 3136
rect 582024 598 582236 626
rect 582024 490 582052 598
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 462 582052 490
rect 582208 480 582236 598
rect 583404 480 583432 3130
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 700304 3478 700360
rect 3054 671200 3110 671256
rect 3238 632032 3294 632088
rect 3330 619112 3386 619168
rect 3238 606056 3294 606112
rect 3146 579944 3202 580000
rect 2870 527856 2926 527912
rect 3238 462576 3294 462632
rect 3330 449520 3386 449576
rect 2962 410488 3018 410544
rect 3238 397432 3294 397488
rect 3330 358400 3386 358456
rect 3146 345344 3202 345400
rect 3330 319232 3386 319288
rect 3054 293120 3110 293176
rect 3146 254088 3202 254144
rect 3054 201864 3110 201920
rect 3514 684256 3570 684312
rect 3514 658180 3516 658200
rect 3516 658180 3568 658200
rect 3568 658180 3570 658200
rect 3514 658144 3570 658180
rect 3514 566888 3570 566944
rect 3514 553832 3570 553888
rect 3514 514800 3570 514856
rect 3514 501744 3570 501800
rect 3514 475632 3570 475688
rect 3514 423580 3516 423600
rect 3516 423580 3568 423600
rect 3568 423580 3570 423600
rect 3514 423544 3570 423580
rect 3514 371320 3570 371376
rect 3514 306176 3570 306232
rect 3514 241032 3570 241088
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 137944 3478 138000
rect 3422 136720 3478 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3330 59200 3386 59256
rect 3330 58520 3386 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3330 33088 3386 33144
rect 3330 32408 3386 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 17222 701528 17278 701584
rect 235446 703704 235502 703760
rect 25502 701664 25558 701720
rect 29642 701392 29698 701448
rect 33782 701256 33838 701312
rect 39394 701120 39450 701176
rect 51722 701800 51778 701856
rect 40498 700984 40554 701040
rect 40682 699760 40738 699816
rect 105450 700712 105506 700768
rect 154118 700848 154174 700904
rect 170310 700576 170366 700632
rect 177302 700168 177358 700224
rect 182730 303456 182786 303512
rect 310886 703568 310942 703624
rect 212630 701936 212686 701992
rect 216126 701936 216182 701992
rect 218978 701936 219034 701992
rect 223118 701936 223174 701992
rect 251178 702480 251234 702536
rect 244002 702344 244058 702400
rect 247682 702344 247738 702400
rect 247866 702344 247922 702400
rect 233606 702072 233662 702128
rect 240690 702072 240746 702128
rect 230110 701936 230166 701992
rect 237194 701936 237250 701992
rect 244186 702208 244242 702264
rect 321374 703432 321430 703488
rect 316130 702480 316186 702536
rect 331862 702888 331918 702944
rect 348974 703432 349030 703488
rect 353298 703432 353354 703488
rect 342442 702752 342498 702808
rect 333978 702616 334034 702672
rect 333242 702480 333298 702536
rect 345938 702480 345994 702536
rect 349066 702480 349122 702536
rect 362958 703024 363014 703080
rect 353114 702752 353170 702808
rect 353298 702752 353354 702808
rect 362222 702616 362278 702672
rect 352930 702480 352986 702536
rect 353114 702480 353170 702536
rect 365718 703840 365774 703896
rect 374642 703840 374698 703896
rect 369674 703024 369730 703080
rect 369490 702616 369546 702672
rect 369674 702616 369730 702672
rect 365810 702480 365866 702536
rect 369674 702500 369730 702536
rect 369674 702480 369676 702500
rect 369676 702480 369728 702500
rect 369728 702480 369730 702500
rect 374090 702480 374146 702536
rect 395066 703704 395122 703760
rect 374642 703024 374698 703080
rect 380990 702480 381046 702536
rect 374642 702344 374698 702400
rect 375378 702344 375434 702400
rect 391110 702480 391166 702536
rect 405554 703432 405610 703488
rect 412638 702616 412694 702672
rect 426622 703296 426678 703352
rect 416134 703160 416190 703216
rect 418066 703160 418122 703216
rect 427634 702616 427690 702672
rect 494794 702752 494850 702808
rect 496910 701664 496966 701720
rect 514114 701800 514170 701856
rect 492954 701528 493010 701584
rect 503626 701528 503682 701584
rect 506938 701392 506994 701448
rect 517610 701392 517666 701448
rect 524602 701256 524658 701312
rect 538954 702208 539010 702264
rect 559654 702480 559710 702536
rect 577042 703468 577044 703488
rect 577044 703468 577096 703488
rect 577096 703468 577098 703488
rect 577042 703432 577098 703468
rect 582470 702072 582526 702128
rect 510710 701120 510766 701176
rect 521106 701120 521162 701176
rect 527178 701120 527234 701176
rect 528190 701120 528246 701176
rect 531962 701120 532018 701176
rect 532238 701156 532240 701176
rect 532240 701156 532292 701176
rect 532292 701156 532294 701176
rect 532238 701120 532294 701156
rect 545578 701120 545634 701176
rect 549718 701120 549774 701176
rect 559838 701120 559894 701176
rect 570234 701120 570290 701176
rect 573730 701120 573786 701176
rect 581090 701120 581146 701176
rect 240874 300192 240930 300248
rect 579802 139340 579804 139360
rect 579804 139340 579856 139360
rect 579856 139340 579858 139360
rect 579802 139304 579858 139340
rect 579986 112784 580042 112840
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 46280 580226 46336
rect 579802 33108 579858 33144
rect 579802 33088 579804 33108
rect 579804 33088 579856 33108
rect 579856 33088 579858 33108
rect 580170 19760 580226 19816
rect 580446 300056 580502 300112
rect 580446 219000 580502 219056
rect 580354 59608 580410 59664
rect 582654 700032 582710 700088
rect 582562 537784 582618 537840
rect 583850 644272 583906 644328
rect 583758 631352 583814 631408
rect 583758 579536 583814 579592
rect 583666 578176 583722 578232
rect 583574 525000 583630 525056
rect 583482 485152 583538 485208
rect 583390 471416 583446 471472
rect 583298 431568 583354 431624
rect 583206 418240 583262 418296
rect 583114 404912 583170 404968
rect 583022 378392 583078 378448
rect 582930 365064 582986 365120
rect 582838 325216 582894 325272
rect 582746 312024 582802 312080
rect 582746 298732 582748 298752
rect 582748 298732 582800 298752
rect 582800 298732 582802 298752
rect 582746 298696 582802 298732
rect 582654 272176 582710 272232
rect 582654 258884 582656 258904
rect 582656 258884 582708 258904
rect 582708 258884 582710 258904
rect 582654 258848 582710 258884
rect 582470 232328 582526 232384
rect 582562 165860 582564 165880
rect 582564 165860 582616 165880
rect 582616 165860 582618 165880
rect 582562 165824 582618 165860
rect 582470 152668 582472 152688
rect 582472 152668 582524 152688
rect 582524 152668 582526 152688
rect 582470 152632 582526 152668
rect 580262 6568 580318 6624
<< metal3 >>
rect 365713 703898 365779 703901
rect 374637 703898 374703 703901
rect 365713 703896 374703 703898
rect 365713 703840 365718 703896
rect 365774 703840 374642 703896
rect 374698 703840 374703 703896
rect 365713 703838 374703 703840
rect 365713 703835 365779 703838
rect 374637 703835 374703 703838
rect 235441 703762 235507 703765
rect 395061 703762 395127 703765
rect 235441 703760 395127 703762
rect 235441 703704 235446 703760
rect 235502 703704 395066 703760
rect 395122 703704 395127 703760
rect 235441 703702 395127 703704
rect 235441 703699 235507 703702
rect 395061 703699 395127 703702
rect 310881 703626 310947 703629
rect 577446 703626 577452 703628
rect 310881 703624 577452 703626
rect 310881 703568 310886 703624
rect 310942 703568 577452 703624
rect 310881 703566 577452 703568
rect 310881 703563 310947 703566
rect 577446 703564 577452 703566
rect 577516 703564 577522 703628
rect 321369 703490 321435 703493
rect 347814 703490 347820 703492
rect 321369 703488 347820 703490
rect 321369 703432 321374 703488
rect 321430 703432 347820 703488
rect 321369 703430 347820 703432
rect 321369 703427 321435 703430
rect 347814 703428 347820 703430
rect 347884 703428 347890 703492
rect 348969 703490 349035 703493
rect 353293 703490 353359 703493
rect 348969 703488 353359 703490
rect 348969 703432 348974 703488
rect 349030 703432 353298 703488
rect 353354 703432 353359 703488
rect 348969 703430 353359 703432
rect 348969 703427 349035 703430
rect 353293 703427 353359 703430
rect 361430 703428 361436 703492
rect 361500 703490 361506 703492
rect 405549 703490 405615 703493
rect 361500 703488 405615 703490
rect 361500 703432 405554 703488
rect 405610 703432 405615 703488
rect 361500 703430 405615 703432
rect 361500 703428 361506 703430
rect 405549 703427 405615 703430
rect 577037 703490 577103 703493
rect 577262 703490 577268 703492
rect 577037 703488 577268 703490
rect 577037 703432 577042 703488
rect 577098 703432 577268 703488
rect 577037 703430 577268 703432
rect 577037 703427 577103 703430
rect 577262 703428 577268 703430
rect 577332 703428 577338 703492
rect 329782 703292 329788 703356
rect 329852 703354 329858 703356
rect 426617 703354 426683 703357
rect 329852 703352 426683 703354
rect 329852 703296 426622 703352
rect 426678 703296 426683 703352
rect 329852 703294 426683 703296
rect 329852 703292 329858 703294
rect 426617 703291 426683 703294
rect 343582 703156 343588 703220
rect 343652 703218 343658 703220
rect 416129 703218 416195 703221
rect 343652 703216 416195 703218
rect 343652 703160 416134 703216
rect 416190 703160 416195 703216
rect 343652 703158 416195 703160
rect 343652 703156 343658 703158
rect 416129 703155 416195 703158
rect 418061 703218 418127 703221
rect 580574 703218 580580 703220
rect 418061 703216 580580 703218
rect 418061 703160 418066 703216
rect 418122 703160 580580 703216
rect 418061 703158 580580 703160
rect 418061 703155 418127 703158
rect 580574 703156 580580 703158
rect 580644 703156 580650 703220
rect 316166 703020 316172 703084
rect 316236 703082 316242 703084
rect 362953 703082 363019 703085
rect 316236 703080 363019 703082
rect 316236 703024 362958 703080
rect 363014 703024 363019 703080
rect 316236 703022 363019 703024
rect 316236 703020 316242 703022
rect 362953 703019 363019 703022
rect 365662 703020 365668 703084
rect 365732 703082 365738 703084
rect 369669 703082 369735 703085
rect 365732 703080 369735 703082
rect 365732 703024 369674 703080
rect 369730 703024 369735 703080
rect 365732 703022 369735 703024
rect 365732 703020 365738 703022
rect 369669 703019 369735 703022
rect 374637 703082 374703 703085
rect 577630 703082 577636 703084
rect 374637 703080 577636 703082
rect 374637 703024 374642 703080
rect 374698 703024 577636 703080
rect 374637 703022 577636 703024
rect 374637 703019 374703 703022
rect 577630 703020 577636 703022
rect 577700 703020 577706 703084
rect 331857 702946 331923 702949
rect 579838 702946 579844 702948
rect 331857 702944 579844 702946
rect 331857 702888 331862 702944
rect 331918 702888 579844 702944
rect 331857 702886 579844 702888
rect 331857 702883 331923 702886
rect 579838 702884 579844 702886
rect 579908 702884 579914 702948
rect 342437 702810 342503 702813
rect 353109 702810 353175 702813
rect 342437 702808 353175 702810
rect 342437 702752 342442 702808
rect 342498 702752 353114 702808
rect 353170 702752 353175 702808
rect 342437 702750 353175 702752
rect 342437 702747 342503 702750
rect 353109 702747 353175 702750
rect 353293 702810 353359 702813
rect 374862 702810 374868 702812
rect 353293 702808 374868 702810
rect 353293 702752 353298 702808
rect 353354 702752 374868 702808
rect 353293 702750 374868 702752
rect 353293 702747 353359 702750
rect 374862 702748 374868 702750
rect 374932 702748 374938 702812
rect 375414 702748 375420 702812
rect 375484 702810 375490 702812
rect 494789 702810 494855 702813
rect 375484 702808 494855 702810
rect 375484 702752 494794 702808
rect 494850 702752 494855 702808
rect 375484 702750 494855 702752
rect 375484 702748 375490 702750
rect 494789 702747 494855 702750
rect 333973 702674 334039 702677
rect 362217 702674 362283 702677
rect 369485 702674 369551 702677
rect 333973 702672 362283 702674
rect 333973 702616 333978 702672
rect 334034 702616 362222 702672
rect 362278 702616 362283 702672
rect 333973 702614 362283 702616
rect 333973 702611 334039 702614
rect 362217 702611 362283 702614
rect 364290 702672 369551 702674
rect 364290 702616 369490 702672
rect 369546 702616 369551 702672
rect 364290 702614 369551 702616
rect 251173 702540 251239 702541
rect 316125 702540 316191 702541
rect 333237 702540 333303 702541
rect 345933 702540 345999 702541
rect 251173 702538 251220 702540
rect 243862 702478 244658 702538
rect 251128 702536 251220 702538
rect 251128 702480 251178 702536
rect 251128 702478 251220 702480
rect 228766 702340 228772 702404
rect 228836 702402 228842 702404
rect 243862 702402 243922 702478
rect 228836 702342 243922 702402
rect 243997 702402 244063 702405
rect 244598 702402 244658 702478
rect 251173 702476 251220 702478
rect 251284 702476 251290 702540
rect 316125 702538 316172 702540
rect 316080 702536 316172 702538
rect 316080 702480 316130 702536
rect 316080 702478 316172 702480
rect 316125 702476 316172 702478
rect 316236 702476 316242 702540
rect 333237 702538 333284 702540
rect 333192 702536 333284 702538
rect 333192 702480 333242 702536
rect 333192 702478 333284 702480
rect 333237 702476 333284 702478
rect 333348 702476 333354 702540
rect 345933 702538 345980 702540
rect 345888 702536 345980 702538
rect 345888 702480 345938 702536
rect 345888 702478 345980 702480
rect 345933 702476 345980 702478
rect 346044 702476 346050 702540
rect 347814 702476 347820 702540
rect 347884 702538 347890 702540
rect 349061 702538 349127 702541
rect 352925 702540 352991 702541
rect 352925 702538 352972 702540
rect 347884 702536 349127 702538
rect 347884 702480 349066 702536
rect 349122 702480 349127 702536
rect 347884 702478 349127 702480
rect 352880 702536 352972 702538
rect 352880 702480 352930 702536
rect 352880 702478 352972 702480
rect 347884 702476 347890 702478
rect 251173 702475 251239 702476
rect 316125 702475 316191 702476
rect 333237 702475 333303 702476
rect 345933 702475 345999 702476
rect 349061 702475 349127 702478
rect 352925 702476 352972 702478
rect 353036 702476 353042 702540
rect 353109 702538 353175 702541
rect 364290 702538 364350 702614
rect 369485 702611 369551 702614
rect 369669 702674 369735 702677
rect 391974 702674 391980 702676
rect 369669 702672 391980 702674
rect 369669 702616 369674 702672
rect 369730 702616 391980 702672
rect 369669 702614 391980 702616
rect 369669 702611 369735 702614
rect 391974 702612 391980 702614
rect 392044 702612 392050 702676
rect 412398 702612 412404 702676
rect 412468 702674 412474 702676
rect 412633 702674 412699 702677
rect 427629 702676 427695 702677
rect 427629 702674 427676 702676
rect 412468 702672 412699 702674
rect 412468 702616 412638 702672
rect 412694 702616 412699 702672
rect 412468 702614 412699 702616
rect 427584 702672 427676 702674
rect 427584 702616 427634 702672
rect 427584 702614 427676 702616
rect 412468 702612 412474 702614
rect 412633 702611 412699 702614
rect 427629 702612 427676 702614
rect 427740 702612 427746 702676
rect 427629 702611 427695 702612
rect 365805 702540 365871 702541
rect 369669 702540 369735 702541
rect 365805 702538 365852 702540
rect 353109 702536 364350 702538
rect 353109 702480 353114 702536
rect 353170 702480 364350 702536
rect 353109 702478 364350 702480
rect 365760 702536 365852 702538
rect 365760 702480 365810 702536
rect 365760 702478 365852 702480
rect 352925 702475 352991 702476
rect 353109 702475 353175 702478
rect 365805 702476 365852 702478
rect 365916 702476 365922 702540
rect 369669 702538 369716 702540
rect 369624 702536 369716 702538
rect 369624 702480 369674 702536
rect 369624 702478 369716 702480
rect 369669 702476 369716 702478
rect 369780 702476 369786 702540
rect 371918 702476 371924 702540
rect 371988 702538 371994 702540
rect 374085 702538 374151 702541
rect 371988 702536 374151 702538
rect 371988 702480 374090 702536
rect 374146 702480 374151 702536
rect 371988 702478 374151 702480
rect 371988 702476 371994 702478
rect 365805 702475 365871 702476
rect 369669 702475 369735 702476
rect 374085 702475 374151 702478
rect 378910 702476 378916 702540
rect 378980 702538 378986 702540
rect 380985 702538 381051 702541
rect 378980 702536 381051 702538
rect 378980 702480 380990 702536
rect 381046 702480 381051 702536
rect 378980 702478 381051 702480
rect 378980 702476 378986 702478
rect 380985 702475 381051 702478
rect 391105 702538 391171 702541
rect 559649 702538 559715 702541
rect 391105 702536 559715 702538
rect 391105 702480 391110 702536
rect 391166 702480 559654 702536
rect 559710 702480 559715 702536
rect 391105 702478 559715 702480
rect 391105 702475 391171 702478
rect 559649 702475 559715 702478
rect 247677 702402 247743 702405
rect 243997 702400 244474 702402
rect 243997 702344 244002 702400
rect 244058 702344 244474 702400
rect 243997 702342 244474 702344
rect 244598 702400 247743 702402
rect 244598 702344 247682 702400
rect 247738 702344 247743 702400
rect 244598 702342 247743 702344
rect 228836 702340 228842 702342
rect 243997 702339 244063 702342
rect 229870 702204 229876 702268
rect 229940 702266 229946 702268
rect 244181 702266 244247 702269
rect 229940 702264 244247 702266
rect 229940 702208 244186 702264
rect 244242 702208 244247 702264
rect 229940 702206 244247 702208
rect 244414 702266 244474 702342
rect 247677 702339 247743 702342
rect 247861 702402 247927 702405
rect 374637 702402 374703 702405
rect 247861 702400 374703 702402
rect 247861 702344 247866 702400
rect 247922 702344 374642 702400
rect 374698 702344 374703 702400
rect 247861 702342 374703 702344
rect 247861 702339 247927 702342
rect 374637 702339 374703 702342
rect 375373 702402 375439 702405
rect 579654 702402 579660 702404
rect 375373 702400 579660 702402
rect 375373 702344 375378 702400
rect 375434 702344 579660 702400
rect 375373 702342 579660 702344
rect 375373 702339 375439 702342
rect 579654 702340 579660 702342
rect 579724 702340 579730 702404
rect 538949 702266 539015 702269
rect 244414 702264 539015 702266
rect 244414 702208 538954 702264
rect 539010 702208 539015 702264
rect 244414 702206 539015 702208
rect 229940 702204 229946 702206
rect 244181 702203 244247 702206
rect 538949 702203 539015 702206
rect 233601 702130 233667 702133
rect 240685 702130 240751 702133
rect 582465 702130 582531 702133
rect 233601 702128 238770 702130
rect 233601 702072 233606 702128
rect 233662 702072 238770 702128
rect 233601 702070 238770 702072
rect 233601 702067 233667 702070
rect 212625 701996 212691 701997
rect 212574 701994 212580 701996
rect 212534 701934 212580 701994
rect 212644 701992 212691 701996
rect 212686 701936 212691 701992
rect 212574 701932 212580 701934
rect 212644 701932 212691 701936
rect 215334 701932 215340 701996
rect 215404 701994 215410 701996
rect 216121 701994 216187 701997
rect 218973 701996 219039 701997
rect 218973 701994 219020 701996
rect 215404 701992 216187 701994
rect 215404 701936 216126 701992
rect 216182 701936 216187 701992
rect 215404 701934 216187 701936
rect 218928 701992 219020 701994
rect 218928 701936 218978 701992
rect 218928 701934 219020 701936
rect 215404 701932 215410 701934
rect 212625 701931 212691 701932
rect 216121 701931 216187 701934
rect 218973 701932 219020 701934
rect 219084 701932 219090 701996
rect 222326 701932 222332 701996
rect 222396 701994 222402 701996
rect 223113 701994 223179 701997
rect 230105 701996 230171 701997
rect 230054 701994 230060 701996
rect 222396 701992 223179 701994
rect 222396 701936 223118 701992
rect 223174 701936 223179 701992
rect 222396 701934 223179 701936
rect 230014 701934 230060 701994
rect 230124 701992 230171 701996
rect 230166 701936 230171 701992
rect 222396 701932 222402 701934
rect 218973 701931 219039 701932
rect 223113 701931 223179 701934
rect 230054 701932 230060 701934
rect 230124 701932 230171 701936
rect 230238 701932 230244 701996
rect 230308 701994 230314 701996
rect 237189 701994 237255 701997
rect 230308 701992 237255 701994
rect 230308 701936 237194 701992
rect 237250 701936 237255 701992
rect 230308 701934 237255 701936
rect 238710 701994 238770 702070
rect 240685 702128 582531 702130
rect 240685 702072 240690 702128
rect 240746 702072 582470 702128
rect 582526 702072 582531 702128
rect 240685 702070 582531 702072
rect 240685 702067 240751 702070
rect 582465 702067 582531 702070
rect 582414 701994 582420 701996
rect 238710 701934 582420 701994
rect 230308 701932 230314 701934
rect 230105 701931 230171 701932
rect 237189 701931 237255 701934
rect 582414 701932 582420 701934
rect 582484 701932 582490 701996
rect 51717 701858 51783 701861
rect 514109 701858 514175 701861
rect 51717 701856 514175 701858
rect 51717 701800 51722 701856
rect 51778 701800 514114 701856
rect 514170 701800 514175 701856
rect 51717 701798 514175 701800
rect 51717 701795 51783 701798
rect 514109 701795 514175 701798
rect 25497 701722 25563 701725
rect 496905 701722 496971 701725
rect 25497 701720 496971 701722
rect 25497 701664 25502 701720
rect 25558 701664 496910 701720
rect 496966 701664 496971 701720
rect 25497 701662 496971 701664
rect 25497 701659 25563 701662
rect 496905 701659 496971 701662
rect 17217 701586 17283 701589
rect 492949 701586 493015 701589
rect 17217 701584 493015 701586
rect 17217 701528 17222 701584
rect 17278 701528 492954 701584
rect 493010 701528 493015 701584
rect 17217 701526 493015 701528
rect 17217 701523 17283 701526
rect 492949 701523 493015 701526
rect 503478 701524 503484 701588
rect 503548 701586 503554 701588
rect 503621 701586 503687 701589
rect 503548 701584 503687 701586
rect 503548 701528 503626 701584
rect 503682 701528 503687 701584
rect 503548 701526 503687 701528
rect 503548 701524 503554 701526
rect 503621 701523 503687 701526
rect 29637 701450 29703 701453
rect 506933 701450 506999 701453
rect 517605 701450 517671 701453
rect 29637 701448 506999 701450
rect 29637 701392 29642 701448
rect 29698 701392 506938 701448
rect 506994 701392 506999 701448
rect 29637 701390 506999 701392
rect 29637 701387 29703 701390
rect 506933 701387 506999 701390
rect 509190 701448 517671 701450
rect 509190 701392 517610 701448
rect 517666 701392 517671 701448
rect 509190 701390 517671 701392
rect 33777 701314 33843 701317
rect 509190 701314 509250 701390
rect 517605 701387 517671 701390
rect 524597 701314 524663 701317
rect 33777 701312 509250 701314
rect 33777 701256 33782 701312
rect 33838 701256 509250 701312
rect 33777 701254 509250 701256
rect 510478 701312 524663 701314
rect 510478 701256 524602 701312
rect 524658 701256 524663 701312
rect 510478 701254 524663 701256
rect 33777 701251 33843 701254
rect 39389 701178 39455 701181
rect 510478 701178 510538 701254
rect 524597 701251 524663 701254
rect 510705 701180 510771 701181
rect 510654 701178 510660 701180
rect 39389 701176 510538 701178
rect 39389 701120 39394 701176
rect 39450 701120 510538 701176
rect 39389 701118 510538 701120
rect 510614 701118 510660 701178
rect 510724 701176 510771 701180
rect 510766 701120 510771 701176
rect 39389 701115 39455 701118
rect 510654 701116 510660 701118
rect 510724 701116 510771 701120
rect 520222 701116 520228 701180
rect 520292 701178 520298 701180
rect 521101 701178 521167 701181
rect 527173 701178 527239 701181
rect 528185 701180 528251 701181
rect 528134 701178 528140 701180
rect 520292 701176 521167 701178
rect 520292 701120 521106 701176
rect 521162 701120 521167 701176
rect 520292 701118 521167 701120
rect 520292 701116 520298 701118
rect 510705 701115 510771 701116
rect 521101 701115 521167 701118
rect 527038 701176 527239 701178
rect 527038 701120 527178 701176
rect 527234 701120 527239 701176
rect 527038 701118 527239 701120
rect 528094 701118 528140 701178
rect 528204 701176 528251 701180
rect 528246 701120 528251 701176
rect 40493 701042 40559 701045
rect 329598 701042 329604 701044
rect 40493 701040 329604 701042
rect 40493 700984 40498 701040
rect 40554 700984 329604 701040
rect 40493 700982 329604 700984
rect 40493 700979 40559 700982
rect 329598 700980 329604 700982
rect 329668 700980 329674 701044
rect 333278 700980 333284 701044
rect 333348 701042 333354 701044
rect 371918 701042 371924 701044
rect 333348 700982 371924 701042
rect 333348 700980 333354 700982
rect 371918 700980 371924 700982
rect 371988 700980 371994 701044
rect 374862 700980 374868 701044
rect 374932 701042 374938 701044
rect 378910 701042 378916 701044
rect 374932 700982 378916 701042
rect 374932 700980 374938 700982
rect 378910 700980 378916 700982
rect 378980 700980 378986 701044
rect 391974 700980 391980 701044
rect 392044 701042 392050 701044
rect 527038 701042 527098 701118
rect 527173 701115 527239 701118
rect 528134 701116 528140 701118
rect 528204 701116 528251 701120
rect 528185 701115 528251 701116
rect 531957 701180 532023 701181
rect 532233 701180 532299 701181
rect 531957 701176 532004 701180
rect 532068 701178 532074 701180
rect 531957 701120 531962 701176
rect 531957 701116 532004 701120
rect 532068 701118 532114 701178
rect 532068 701116 532074 701118
rect 532182 701116 532188 701180
rect 532252 701178 532299 701180
rect 532252 701176 532344 701178
rect 532294 701120 532344 701176
rect 532252 701118 532344 701120
rect 532252 701116 532299 701118
rect 545062 701116 545068 701180
rect 545132 701178 545138 701180
rect 545573 701178 545639 701181
rect 545132 701176 545639 701178
rect 545132 701120 545578 701176
rect 545634 701120 545639 701176
rect 545132 701118 545639 701120
rect 545132 701116 545138 701118
rect 531957 701115 532023 701116
rect 532233 701115 532299 701116
rect 545573 701115 545639 701118
rect 549713 701178 549779 701181
rect 559833 701180 559899 701181
rect 550030 701178 550036 701180
rect 549713 701176 550036 701178
rect 549713 701120 549718 701176
rect 549774 701120 550036 701176
rect 549713 701118 550036 701120
rect 549713 701115 549779 701118
rect 550030 701116 550036 701118
rect 550100 701116 550106 701180
rect 559782 701178 559788 701180
rect 559742 701118 559788 701178
rect 559852 701176 559899 701180
rect 559894 701120 559899 701176
rect 559782 701116 559788 701118
rect 559852 701116 559899 701120
rect 570086 701116 570092 701180
rect 570156 701178 570162 701180
rect 570229 701178 570295 701181
rect 570156 701176 570295 701178
rect 570156 701120 570234 701176
rect 570290 701120 570295 701176
rect 570156 701118 570295 701120
rect 570156 701116 570162 701118
rect 559833 701115 559899 701116
rect 570229 701115 570295 701118
rect 572662 701116 572668 701180
rect 572732 701178 572738 701180
rect 573725 701178 573791 701181
rect 572732 701176 573791 701178
rect 572732 701120 573730 701176
rect 573786 701120 573791 701176
rect 572732 701118 573791 701120
rect 572732 701116 572738 701118
rect 573725 701115 573791 701118
rect 580942 701116 580948 701180
rect 581012 701178 581018 701180
rect 581085 701178 581151 701181
rect 581012 701176 581151 701178
rect 581012 701120 581090 701176
rect 581146 701120 581151 701176
rect 581012 701118 581151 701120
rect 581012 701116 581018 701118
rect 581085 701115 581151 701118
rect 392044 700982 527098 701042
rect 392044 700980 392050 700982
rect 154113 700906 154179 700909
rect 412398 700906 412404 700908
rect 154113 700904 412404 700906
rect 154113 700848 154118 700904
rect 154174 700848 412404 700904
rect 154113 700846 412404 700848
rect 154113 700843 154179 700846
rect 412398 700844 412404 700846
rect 412468 700844 412474 700908
rect 427670 700844 427676 700908
rect 427740 700906 427746 700908
rect 580022 700906 580028 700908
rect 427740 700846 580028 700906
rect 427740 700844 427746 700846
rect 580022 700844 580028 700846
rect 580092 700844 580098 700908
rect 105445 700770 105511 700773
rect 343582 700770 343588 700772
rect 105445 700768 343588 700770
rect 105445 700712 105450 700768
rect 105506 700712 343588 700768
rect 105445 700710 343588 700712
rect 105445 700707 105511 700710
rect 343582 700708 343588 700710
rect 343652 700708 343658 700772
rect 345974 700708 345980 700772
rect 346044 700770 346050 700772
rect 365662 700770 365668 700772
rect 346044 700710 365668 700770
rect 346044 700708 346050 700710
rect 365662 700708 365668 700710
rect 365732 700708 365738 700772
rect 369710 700708 369716 700772
rect 369780 700770 369786 700772
rect 580390 700770 580396 700772
rect 369780 700710 580396 700770
rect 369780 700708 369786 700710
rect 580390 700708 580396 700710
rect 580460 700708 580466 700772
rect 170305 700634 170371 700637
rect 361430 700634 361436 700636
rect 170305 700632 361436 700634
rect 170305 700576 170310 700632
rect 170366 700576 361436 700632
rect 170305 700574 361436 700576
rect 170305 700571 170371 700574
rect 361430 700572 361436 700574
rect 361500 700572 361506 700636
rect 365846 700572 365852 700636
rect 365916 700634 365922 700636
rect 580206 700634 580212 700636
rect 365916 700574 580212 700634
rect 365916 700572 365922 700574
rect 580206 700572 580212 700574
rect 580276 700572 580282 700636
rect 219014 700436 219020 700500
rect 219084 700498 219090 700500
rect 315798 700498 315804 700500
rect 219084 700438 315804 700498
rect 219084 700436 219090 700438
rect 315798 700436 315804 700438
rect 315868 700436 315874 700500
rect 316166 700436 316172 700500
rect 316236 700498 316242 700500
rect 559782 700498 559788 700500
rect 316236 700438 559788 700498
rect 316236 700436 316242 700438
rect 559782 700436 559788 700438
rect 559852 700436 559858 700500
rect 3417 700362 3483 700365
rect 532182 700362 532188 700364
rect 3417 700360 532188 700362
rect 3417 700304 3422 700360
rect 3478 700304 532188 700360
rect 3417 700302 532188 700304
rect 3417 700299 3483 700302
rect 532182 700300 532188 700302
rect 532252 700300 532258 700364
rect 177297 700226 177363 700229
rect 503478 700226 503484 700228
rect 177297 700224 503484 700226
rect 177297 700168 177302 700224
rect 177358 700168 503484 700224
rect 177297 700166 503484 700168
rect 177297 700163 177363 700166
rect 503478 700164 503484 700166
rect 503548 700164 503554 700228
rect 251214 700028 251220 700092
rect 251284 700090 251290 700092
rect 582649 700090 582715 700093
rect 251284 700088 582715 700090
rect 251284 700032 582654 700088
rect 582710 700032 582715 700088
rect 251284 700030 582715 700032
rect 251284 700028 251290 700030
rect 582649 700027 582715 700030
rect 230054 699892 230060 699956
rect 230124 699954 230130 699956
rect 582598 699954 582604 699956
rect 230124 699894 582604 699954
rect 230124 699892 230130 699894
rect 582598 699892 582604 699894
rect 582668 699892 582674 699956
rect 40677 699818 40743 699821
rect 528134 699818 528140 699820
rect 40677 699816 528140 699818
rect 40677 699760 40682 699816
rect 40738 699760 528140 699816
rect 40677 699758 528140 699760
rect 40677 699755 40743 699758
rect 528134 699756 528140 699758
rect 528204 699756 528210 699820
rect 352966 699620 352972 699684
rect 353036 699682 353042 699684
rect 375414 699682 375420 699684
rect 353036 699622 375420 699682
rect 353036 699620 353042 699622
rect 375414 699620 375420 699622
rect 375484 699620 375490 699684
rect 579838 697580 579844 697644
rect 579908 697642 579914 697644
rect 580758 697642 580764 697644
rect 579908 697582 580764 697642
rect 579908 697580 579914 697582
rect 580758 697580 580764 697582
rect 580828 697580 580834 697644
rect -960 697220 480 697460
rect 580206 697172 580212 697236
rect 580276 697234 580282 697236
rect 583520 697234 584960 697324
rect 580276 697174 584960 697234
rect 580276 697172 580282 697174
rect 583520 697084 584960 697174
rect 579654 696492 579660 696556
rect 579724 696554 579730 696556
rect 580390 696554 580396 696556
rect 579724 696494 580396 696554
rect 579724 696492 579730 696494
rect 580390 696492 580396 696494
rect 580460 696492 580466 696556
rect -960 684314 480 684404
rect 3509 684314 3575 684317
rect -960 684312 3575 684314
rect -960 684256 3514 684312
rect 3570 684256 3575 684312
rect -960 684254 3575 684256
rect -960 684164 480 684254
rect 3509 684251 3575 684254
rect 580022 683844 580028 683908
rect 580092 683906 580098 683908
rect 583520 683906 584960 683996
rect 580092 683846 584960 683906
rect 580092 683844 580098 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3049 671258 3115 671261
rect -960 671256 3115 671258
rect -960 671200 3054 671256
rect 3110 671200 3115 671256
rect -960 671198 3115 671200
rect -960 671108 480 671198
rect 3049 671195 3115 671198
rect 580758 670652 580764 670716
rect 580828 670714 580834 670716
rect 583520 670714 584960 670804
rect 580828 670654 584960 670714
rect 580828 670652 580834 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583845 644330 583911 644333
rect 583710 644328 583911 644330
rect 583710 644272 583850 644328
rect 583906 644272 583911 644328
rect 583710 644270 583911 644272
rect 583710 644194 583770 644270
rect 583845 644267 583911 644270
rect 583342 644148 583770 644194
rect 583342 644134 584960 644148
rect 583342 644058 583402 644134
rect 583520 644058 584960 644134
rect 583342 643998 584960 644058
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3233 632090 3299 632093
rect -960 632088 3299 632090
rect -960 632032 3238 632088
rect 3294 632032 3299 632088
rect -960 632030 3299 632032
rect -960 631940 480 632030
rect 3233 632027 3299 632030
rect 583753 631410 583819 631413
rect 583710 631408 583819 631410
rect 583710 631352 583758 631408
rect 583814 631352 583819 631408
rect 583710 631347 583819 631352
rect 583710 631002 583770 631347
rect 583342 630956 583770 631002
rect 583342 630942 584960 630956
rect 583342 630866 583402 630942
rect 583520 630866 584960 630942
rect 583342 630806 584960 630866
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3325 619170 3391 619173
rect -960 619168 3391 619170
rect -960 619112 3330 619168
rect 3386 619112 3391 619168
rect -960 619110 3391 619112
rect -960 619020 480 619110
rect 3325 619107 3391 619110
rect 577998 617476 578004 617540
rect 578068 617538 578074 617540
rect 583520 617538 584960 617628
rect 578068 617478 584960 617538
rect 578068 617476 578074 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580574 590956 580580 591020
rect 580644 591018 580650 591020
rect 583520 591018 584960 591108
rect 580644 590958 584960 591018
rect 580644 590956 580650 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3141 580002 3207 580005
rect -960 580000 3207 580002
rect -960 579944 3146 580000
rect 3202 579944 3207 580000
rect -960 579942 3207 579944
rect -960 579852 480 579942
rect 3141 579939 3207 579942
rect 580942 579532 580948 579596
rect 581012 579594 581018 579596
rect 583753 579594 583819 579597
rect 581012 579592 583819 579594
rect 581012 579536 583758 579592
rect 583814 579536 583819 579592
rect 581012 579534 583819 579536
rect 581012 579532 581018 579534
rect 583753 579531 583819 579534
rect 583661 578234 583727 578237
rect 583526 578232 583727 578234
rect 583526 578176 583666 578232
rect 583722 578176 583727 578232
rect 583526 578174 583727 578176
rect 583526 577826 583586 578174
rect 583661 578171 583727 578174
rect 583342 577780 583586 577826
rect 583342 577766 584960 577780
rect 583342 577690 583402 577766
rect 583520 577690 584960 577766
rect 583342 577630 584960 577690
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 577998 564300 578004 564364
rect 578068 564362 578074 564364
rect 583520 564362 584960 564452
rect 578068 564302 584960 564362
rect 578068 564300 578074 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3509 553890 3575 553893
rect -960 553888 3575 553890
rect -960 553832 3514 553888
rect 3570 553832 3575 553888
rect -960 553830 3575 553832
rect -960 553740 480 553830
rect 3509 553827 3575 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 582557 537842 582623 537845
rect 583520 537842 584960 537932
rect 582557 537840 584960 537842
rect 582557 537784 582562 537840
rect 582618 537784 584960 537840
rect 582557 537782 584960 537784
rect 582557 537779 582623 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2865 527914 2931 527917
rect -960 527912 2931 527914
rect -960 527856 2870 527912
rect 2926 527856 2931 527912
rect -960 527854 2931 527856
rect -960 527764 480 527854
rect 2865 527851 2931 527854
rect 583569 525058 583635 525061
rect 583526 525056 583635 525058
rect 583526 525000 583574 525056
rect 583630 525000 583635 525056
rect 583526 524995 583635 525000
rect 583526 524650 583586 524995
rect 583342 524604 583586 524650
rect 583342 524590 584960 524604
rect 583342 524514 583402 524590
rect 583520 524514 584960 524590
rect 583342 524454 584960 524514
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580390 511260 580396 511324
rect 580460 511322 580466 511324
rect 583520 511322 584960 511412
rect 580460 511262 584960 511322
rect 580460 511260 580466 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583477 485210 583543 485213
rect 583477 485208 583586 485210
rect 583477 485152 583482 485208
rect 583538 485152 583586 485208
rect 583477 485147 583586 485152
rect 583526 484802 583586 485147
rect 583342 484756 583586 484802
rect 583342 484742 584960 484756
rect 583342 484666 583402 484742
rect 583520 484666 584960 484742
rect 583342 484606 584960 484666
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3509 475690 3575 475693
rect -960 475688 3575 475690
rect -960 475632 3514 475688
rect 3570 475632 3575 475688
rect -960 475630 3575 475632
rect -960 475540 480 475630
rect 3509 475627 3575 475630
rect 583385 471474 583451 471477
rect 583520 471474 584960 471564
rect 583385 471472 584960 471474
rect 583385 471416 583390 471472
rect 583446 471416 584960 471472
rect 583385 471414 584960 471416
rect 583385 471411 583451 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580206 458084 580212 458148
rect 580276 458146 580282 458148
rect 583520 458146 584960 458236
rect 580276 458086 584960 458146
rect 580276 458084 580282 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583293 431626 583359 431629
rect 583520 431626 584960 431716
rect 583293 431624 584960 431626
rect 583293 431568 583298 431624
rect 583354 431568 584960 431624
rect 583293 431566 584960 431568
rect 583293 431563 583359 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 583201 418298 583267 418301
rect 583520 418298 584960 418388
rect 583201 418296 584960 418298
rect 583201 418240 583206 418296
rect 583262 418240 584960 418296
rect 583201 418238 584960 418240
rect 583201 418235 583267 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 583109 404970 583175 404973
rect 583520 404970 584960 405060
rect 583109 404968 584960 404970
rect 583109 404912 583114 404968
rect 583170 404912 584960 404968
rect 583109 404910 584960 404912
rect 583109 404907 583175 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3233 397490 3299 397493
rect -960 397488 3299 397490
rect -960 397432 3238 397488
rect 3294 397432 3299 397488
rect -960 397430 3299 397432
rect -960 397340 480 397430
rect 3233 397427 3299 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583017 378450 583083 378453
rect 583520 378450 584960 378540
rect 583017 378448 584960 378450
rect 583017 378392 583022 378448
rect 583078 378392 584960 378448
rect 583017 378390 584960 378392
rect 583017 378387 583083 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 582925 365122 582991 365125
rect 583520 365122 584960 365212
rect 582925 365120 584960 365122
rect 582925 365064 582930 365120
rect 582986 365064 584960 365120
rect 582925 365062 584960 365064
rect 582925 365059 582991 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 577998 351868 578004 351932
rect 578068 351930 578074 351932
rect 583520 351930 584960 352020
rect 578068 351870 584960 351930
rect 578068 351868 578074 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 582833 325274 582899 325277
rect 583520 325274 584960 325364
rect 582833 325272 584960 325274
rect 582833 325216 582838 325272
rect 582894 325216 584960 325272
rect 582833 325214 584960 325216
rect 582833 325211 582899 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 582741 312082 582807 312085
rect 583520 312082 584960 312172
rect 582741 312080 584960 312082
rect 582741 312024 582746 312080
rect 582802 312024 584960 312080
rect 582741 312022 584960 312024
rect 582741 312019 582807 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 182725 303514 182791 303517
rect 510654 303514 510660 303516
rect 182725 303512 510660 303514
rect 182725 303456 182730 303512
rect 182786 303456 510660 303512
rect 182725 303454 510660 303456
rect 182725 303451 182791 303454
rect 510654 303452 510660 303454
rect 510724 303452 510730 303516
rect 222326 300188 222332 300252
rect 222396 300250 222402 300252
rect 240869 300250 240935 300253
rect 222396 300248 240935 300250
rect 222396 300192 240874 300248
rect 240930 300192 240935 300248
rect 222396 300190 240935 300192
rect 222396 300188 222402 300190
rect 240869 300187 240935 300190
rect 230054 300052 230060 300116
rect 230124 300114 230130 300116
rect 580441 300114 580507 300117
rect 230124 300112 580507 300114
rect 230124 300056 580446 300112
rect 580502 300056 580507 300112
rect 230124 300054 580507 300056
rect 230124 300052 230130 300054
rect 580441 300051 580507 300054
rect 582741 298754 582807 298757
rect 583520 298754 584960 298844
rect 582741 298752 584960 298754
rect 582741 298696 582746 298752
rect 582802 298696 584960 298752
rect 582741 298694 584960 298696
rect 582741 298691 582807 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 582649 272234 582715 272237
rect 583520 272234 584960 272324
rect 582649 272232 584960 272234
rect 582649 272176 582654 272232
rect 582710 272176 584960 272232
rect 582649 272174 584960 272176
rect 582649 272171 582715 272174
rect 583520 272084 584960 272174
rect 520222 267746 520228 267748
rect 430 267686 520228 267746
rect 430 267474 490 267686
rect 520222 267684 520228 267686
rect 520292 267684 520298 267748
rect 430 267414 674 267474
rect -960 267202 480 267292
rect 614 267202 674 267414
rect -960 267142 674 267202
rect -960 267052 480 267142
rect 582649 258906 582715 258909
rect 583520 258906 584960 258996
rect 582649 258904 584960 258906
rect 582649 258848 582654 258904
rect 582710 258848 584960 258904
rect 582649 258846 584960 258848
rect 582649 258843 582715 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 583520 245578 584960 245668
rect 583342 245518 584960 245578
rect 583342 245442 583402 245518
rect 583520 245442 584960 245518
rect 583342 245428 584960 245442
rect 583342 245382 583586 245428
rect 228766 244292 228772 244356
rect 228836 244354 228842 244356
rect 583526 244354 583586 245382
rect 228836 244294 583586 244354
rect 228836 244292 228842 244294
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 582465 232386 582531 232389
rect 583520 232386 584960 232476
rect 582465 232384 584960 232386
rect 582465 232328 582470 232384
rect 582526 232328 584960 232384
rect 582465 232326 584960 232328
rect 582465 232323 582531 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580441 219058 580507 219061
rect 583520 219058 584960 219148
rect 580441 219056 584960 219058
rect 580441 219000 580446 219056
rect 580502 219000 584960 219056
rect 580441 218998 584960 219000
rect 580441 218995 580507 218998
rect 583520 218908 584960 218998
rect 531998 215250 532004 215252
rect 6870 215190 532004 215250
rect -960 214978 480 215068
rect 6870 214978 6930 215190
rect 531998 215188 532004 215190
rect 532068 215188 532074 215252
rect -960 214918 6930 214978
rect -960 214828 480 214918
rect 230238 205668 230244 205732
rect 230308 205730 230314 205732
rect 583520 205730 584960 205820
rect 230308 205670 584960 205730
rect 230308 205668 230314 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 582598 192476 582604 192540
rect 582668 192538 582674 192540
rect 583520 192538 584960 192628
rect 582668 192478 584960 192538
rect 582668 192476 582674 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 582414 179148 582420 179212
rect 582484 179210 582490 179212
rect 583520 179210 584960 179300
rect 582484 179150 584960 179210
rect 582484 179148 582490 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 582557 165882 582623 165885
rect 583520 165882 584960 165972
rect 582557 165880 584960 165882
rect 582557 165824 582562 165880
rect 582618 165824 584960 165880
rect 582557 165822 584960 165824
rect 582557 165819 582623 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 582465 152690 582531 152693
rect 583520 152690 584960 152780
rect 582465 152688 584960 152690
rect 582465 152632 582470 152688
rect 582526 152632 584960 152688
rect 582465 152630 584960 152632
rect 582465 152627 582531 152630
rect 583520 152540 584960 152630
rect 550030 150378 550036 150380
rect 430 150318 550036 150378
rect 430 150106 490 150318
rect 550030 150316 550036 150318
rect 550100 150316 550106 150380
rect 430 150046 674 150106
rect -960 149834 480 149924
rect 614 149834 674 150046
rect -960 149774 674 149834
rect -960 149684 480 149774
rect 579797 139362 579863 139365
rect 583520 139362 584960 139452
rect 579797 139360 584960 139362
rect 579797 139304 579802 139360
rect 579858 139304 584960 139360
rect 579797 139302 584960 139304
rect 579797 139299 579863 139302
rect 583520 139212 584960 139302
rect 3417 138002 3483 138005
rect 545062 138002 545068 138004
rect 3417 138000 545068 138002
rect 3417 137944 3422 138000
rect 3478 137944 545068 138000
rect 3417 137942 545068 137944
rect 3417 137939 3483 137942
rect 545062 137940 545068 137942
rect 545132 137940 545138 138004
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 583520 126034 584960 126124
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 215334 125564 215340 125628
rect 215404 125626 215410 125628
rect 583526 125626 583586 125838
rect 215404 125566 583586 125626
rect 215404 125564 215410 125566
rect -960 123572 480 123812
rect 579981 112842 580047 112845
rect 583520 112842 584960 112932
rect 579981 112840 584960 112842
rect 579981 112784 579986 112840
rect 580042 112784 584960 112840
rect 579981 112782 584960 112784
rect 579981 112779 580047 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 212574 99452 212580 99516
rect 212644 99514 212650 99516
rect 583520 99514 584960 99604
rect 212644 99454 584960 99514
rect 212644 99452 212650 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580349 59666 580415 59669
rect 583520 59666 584960 59756
rect 580349 59664 584960 59666
rect 580349 59608 580354 59664
rect 580410 59608 584960 59664
rect 580349 59606 584960 59608
rect 580349 59603 580415 59606
rect 583520 59516 584960 59606
rect 3325 59258 3391 59261
rect 570086 59258 570092 59260
rect 3325 59256 570092 59258
rect 3325 59200 3330 59256
rect 3386 59200 570092 59256
rect 3325 59198 570092 59200
rect 3325 59195 3391 59198
rect 570086 59196 570092 59198
rect 570156 59196 570162 59260
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 3325 33146 3391 33149
rect 572662 33146 572668 33148
rect 3325 33144 572668 33146
rect 3325 33088 3330 33144
rect 3386 33088 572668 33144
rect 3325 33086 572668 33088
rect 3325 33083 3391 33086
rect 572662 33084 572668 33086
rect 572732 33084 572738 33148
rect 579797 33146 579863 33149
rect 583520 33146 584960 33236
rect 579797 33144 584960 33146
rect 579797 33088 579802 33144
rect 579858 33088 584960 33144
rect 579797 33086 584960 33088
rect 579797 33083 579863 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3325 32466 3391 32469
rect -960 32464 3391 32466
rect -960 32408 3330 32464
rect 3386 32408 3391 32464
rect -960 32406 3391 32408
rect -960 32316 480 32406
rect 3325 32403 3391 32406
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 577452 703564 577516 703628
rect 347820 703428 347884 703492
rect 361436 703428 361500 703492
rect 577268 703428 577332 703492
rect 329788 703292 329852 703356
rect 343588 703156 343652 703220
rect 580580 703156 580644 703220
rect 316172 703020 316236 703084
rect 365668 703020 365732 703084
rect 577636 703020 577700 703084
rect 579844 702884 579908 702948
rect 374868 702748 374932 702812
rect 375420 702748 375484 702812
rect 251220 702536 251284 702540
rect 251220 702480 251234 702536
rect 251234 702480 251284 702536
rect 228772 702340 228836 702404
rect 251220 702476 251284 702480
rect 316172 702536 316236 702540
rect 316172 702480 316186 702536
rect 316186 702480 316236 702536
rect 316172 702476 316236 702480
rect 333284 702536 333348 702540
rect 333284 702480 333298 702536
rect 333298 702480 333348 702536
rect 333284 702476 333348 702480
rect 345980 702536 346044 702540
rect 345980 702480 345994 702536
rect 345994 702480 346044 702536
rect 345980 702476 346044 702480
rect 347820 702476 347884 702540
rect 352972 702536 353036 702540
rect 352972 702480 352986 702536
rect 352986 702480 353036 702536
rect 352972 702476 353036 702480
rect 391980 702612 392044 702676
rect 412404 702612 412468 702676
rect 427676 702672 427740 702676
rect 427676 702616 427690 702672
rect 427690 702616 427740 702672
rect 427676 702612 427740 702616
rect 365852 702536 365916 702540
rect 365852 702480 365866 702536
rect 365866 702480 365916 702536
rect 365852 702476 365916 702480
rect 369716 702536 369780 702540
rect 369716 702480 369730 702536
rect 369730 702480 369780 702536
rect 369716 702476 369780 702480
rect 371924 702476 371988 702540
rect 378916 702476 378980 702540
rect 229876 702204 229940 702268
rect 579660 702340 579724 702404
rect 212580 701992 212644 701996
rect 212580 701936 212630 701992
rect 212630 701936 212644 701992
rect 212580 701932 212644 701936
rect 215340 701932 215404 701996
rect 219020 701992 219084 701996
rect 219020 701936 219034 701992
rect 219034 701936 219084 701992
rect 219020 701932 219084 701936
rect 222332 701932 222396 701996
rect 230060 701992 230124 701996
rect 230060 701936 230110 701992
rect 230110 701936 230124 701992
rect 230060 701932 230124 701936
rect 230244 701932 230308 701996
rect 582420 701932 582484 701996
rect 503484 701524 503548 701588
rect 510660 701176 510724 701180
rect 510660 701120 510710 701176
rect 510710 701120 510724 701176
rect 510660 701116 510724 701120
rect 520228 701116 520292 701180
rect 528140 701176 528204 701180
rect 528140 701120 528190 701176
rect 528190 701120 528204 701176
rect 329604 700980 329668 701044
rect 333284 700980 333348 701044
rect 371924 700980 371988 701044
rect 374868 700980 374932 701044
rect 378916 700980 378980 701044
rect 391980 700980 392044 701044
rect 528140 701116 528204 701120
rect 532004 701176 532068 701180
rect 532004 701120 532018 701176
rect 532018 701120 532068 701176
rect 532004 701116 532068 701120
rect 532188 701176 532252 701180
rect 532188 701120 532238 701176
rect 532238 701120 532252 701176
rect 532188 701116 532252 701120
rect 545068 701116 545132 701180
rect 550036 701116 550100 701180
rect 559788 701176 559852 701180
rect 559788 701120 559838 701176
rect 559838 701120 559852 701176
rect 559788 701116 559852 701120
rect 570092 701116 570156 701180
rect 572668 701116 572732 701180
rect 580948 701116 581012 701180
rect 412404 700844 412468 700908
rect 427676 700844 427740 700908
rect 580028 700844 580092 700908
rect 343588 700708 343652 700772
rect 345980 700708 346044 700772
rect 365668 700708 365732 700772
rect 369716 700708 369780 700772
rect 580396 700708 580460 700772
rect 361436 700572 361500 700636
rect 365852 700572 365916 700636
rect 580212 700572 580276 700636
rect 219020 700436 219084 700500
rect 315804 700436 315868 700500
rect 316172 700436 316236 700500
rect 559788 700436 559852 700500
rect 532188 700300 532252 700364
rect 503484 700164 503548 700228
rect 251220 700028 251284 700092
rect 230060 699892 230124 699956
rect 582604 699892 582668 699956
rect 528140 699756 528204 699820
rect 352972 699620 353036 699684
rect 375420 699620 375484 699684
rect 579844 697580 579908 697644
rect 580764 697580 580828 697644
rect 580212 697172 580276 697236
rect 579660 696492 579724 696556
rect 580396 696492 580460 696556
rect 580028 683844 580092 683908
rect 580764 670652 580828 670716
rect 578004 617476 578068 617540
rect 580580 590956 580644 591020
rect 580948 579532 581012 579596
rect 578004 564300 578068 564364
rect 580396 511260 580460 511324
rect 580212 458084 580276 458148
rect 578004 351868 578068 351932
rect 510660 303452 510724 303516
rect 222332 300188 222396 300252
rect 230060 300052 230124 300116
rect 520228 267684 520292 267748
rect 228772 244292 228836 244356
rect 532004 215188 532068 215252
rect 230244 205668 230308 205732
rect 582604 192476 582668 192540
rect 582420 179148 582484 179212
rect 550036 150316 550100 150380
rect 545068 137940 545132 138004
rect 215340 125564 215404 125628
rect 212580 99452 212644 99516
rect 570092 59196 570156 59260
rect 572668 33084 572732 33148
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 185514 703784 186134 706202
rect 189234 703784 189854 708122
rect 192954 703784 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 701784 200414 705242
rect 203514 703784 204134 707162
rect 207234 703784 207854 709082
rect 210954 703784 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 212579 701996 212645 701997
rect 212579 701932 212580 701996
rect 212644 701932 212645 701996
rect 212579 701931 212645 701932
rect 215339 701996 215405 701997
rect 215339 701932 215340 701996
rect 215404 701932 215405 701996
rect 215339 701931 215405 701932
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 186992 687454 187312 687486
rect 186992 687218 187034 687454
rect 187270 687218 187312 687454
rect 186992 687134 187312 687218
rect 186992 686898 187034 687134
rect 187270 686898 187312 687134
rect 186992 686866 187312 686898
rect 202352 669454 202672 669486
rect 202352 669218 202394 669454
rect 202630 669218 202672 669454
rect 202352 669134 202672 669218
rect 202352 668898 202394 669134
rect 202630 668898 202672 669134
rect 202352 668866 202672 668898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 186992 651454 187312 651486
rect 186992 651218 187034 651454
rect 187270 651218 187312 651454
rect 186992 651134 187312 651218
rect 186992 650898 187034 651134
rect 187270 650898 187312 651134
rect 186992 650866 187312 650898
rect 202352 633454 202672 633486
rect 202352 633218 202394 633454
rect 202630 633218 202672 633454
rect 202352 633134 202672 633218
rect 202352 632898 202394 633134
rect 202630 632898 202672 633134
rect 202352 632866 202672 632898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 186992 615454 187312 615486
rect 186992 615218 187034 615454
rect 187270 615218 187312 615454
rect 186992 615134 187312 615218
rect 186992 614898 187034 615134
rect 187270 614898 187312 615134
rect 186992 614866 187312 614898
rect 202352 597454 202672 597486
rect 202352 597218 202394 597454
rect 202630 597218 202672 597454
rect 202352 597134 202672 597218
rect 202352 596898 202394 597134
rect 202630 596898 202672 597134
rect 202352 596866 202672 596898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 186992 579454 187312 579486
rect 186992 579218 187034 579454
rect 187270 579218 187312 579454
rect 186992 579134 187312 579218
rect 186992 578898 187034 579134
rect 187270 578898 187312 579134
rect 186992 578866 187312 578898
rect 202352 561454 202672 561486
rect 202352 561218 202394 561454
rect 202630 561218 202672 561454
rect 202352 561134 202672 561218
rect 202352 560898 202394 561134
rect 202630 560898 202672 561134
rect 202352 560866 202672 560898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 186992 543454 187312 543486
rect 186992 543218 187034 543454
rect 187270 543218 187312 543454
rect 186992 543134 187312 543218
rect 186992 542898 187034 543134
rect 187270 542898 187312 543134
rect 186992 542866 187312 542898
rect 202352 525454 202672 525486
rect 202352 525218 202394 525454
rect 202630 525218 202672 525454
rect 202352 525134 202672 525218
rect 202352 524898 202394 525134
rect 202630 524898 202672 525134
rect 202352 524866 202672 524898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 186992 507454 187312 507486
rect 186992 507218 187034 507454
rect 187270 507218 187312 507454
rect 186992 507134 187312 507218
rect 186992 506898 187034 507134
rect 187270 506898 187312 507134
rect 186992 506866 187312 506898
rect 202352 489454 202672 489486
rect 202352 489218 202394 489454
rect 202630 489218 202672 489454
rect 202352 489134 202672 489218
rect 202352 488898 202394 489134
rect 202630 488898 202672 489134
rect 202352 488866 202672 488898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 186992 471454 187312 471486
rect 186992 471218 187034 471454
rect 187270 471218 187312 471454
rect 186992 471134 187312 471218
rect 186992 470898 187034 471134
rect 187270 470898 187312 471134
rect 186992 470866 187312 470898
rect 202352 453454 202672 453486
rect 202352 453218 202394 453454
rect 202630 453218 202672 453454
rect 202352 453134 202672 453218
rect 202352 452898 202394 453134
rect 202630 452898 202672 453134
rect 202352 452866 202672 452898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 186992 435454 187312 435486
rect 186992 435218 187034 435454
rect 187270 435218 187312 435454
rect 186992 435134 187312 435218
rect 186992 434898 187034 435134
rect 187270 434898 187312 435134
rect 186992 434866 187312 434898
rect 202352 417454 202672 417486
rect 202352 417218 202394 417454
rect 202630 417218 202672 417454
rect 202352 417134 202672 417218
rect 202352 416898 202394 417134
rect 202630 416898 202672 417134
rect 202352 416866 202672 416898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 186992 399454 187312 399486
rect 186992 399218 187034 399454
rect 187270 399218 187312 399454
rect 186992 399134 187312 399218
rect 186992 398898 187034 399134
rect 187270 398898 187312 399134
rect 186992 398866 187312 398898
rect 202352 381454 202672 381486
rect 202352 381218 202394 381454
rect 202630 381218 202672 381454
rect 202352 381134 202672 381218
rect 202352 380898 202394 381134
rect 202630 380898 202672 381134
rect 202352 380866 202672 380898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 186992 363454 187312 363486
rect 186992 363218 187034 363454
rect 187270 363218 187312 363454
rect 186992 363134 187312 363218
rect 186992 362898 187034 363134
rect 187270 362898 187312 363134
rect 186992 362866 187312 362898
rect 202352 345454 202672 345486
rect 202352 345218 202394 345454
rect 202630 345218 202672 345454
rect 202352 345134 202672 345218
rect 202352 344898 202394 345134
rect 202630 344898 202672 345134
rect 202352 344866 202672 344898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 186992 327454 187312 327486
rect 186992 327218 187034 327454
rect 187270 327218 187312 327454
rect 186992 327134 187312 327218
rect 186992 326898 187034 327134
rect 187270 326898 187312 327134
rect 186992 326866 187312 326898
rect 202352 309454 202672 309486
rect 202352 309218 202394 309454
rect 202630 309218 202672 309454
rect 202352 309134 202672 309218
rect 202352 308898 202394 309134
rect 202630 308898 202672 309134
rect 202352 308866 202672 308898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 295174 186134 299784
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 298894 189854 299784
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 266614 193574 299784
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 273454 200414 301784
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 277174 204134 299784
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 280894 207854 299784
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 284614 211574 299784
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 212582 99517 212642 701931
rect 215342 125629 215402 701931
rect 217794 701784 218414 704282
rect 221514 703784 222134 706202
rect 225234 703784 225854 708122
rect 228954 703784 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 228771 702404 228837 702405
rect 228771 702340 228772 702404
rect 228836 702340 228837 702404
rect 228771 702339 228837 702340
rect 219019 701996 219085 701997
rect 219019 701932 219020 701996
rect 219084 701932 219085 701996
rect 219019 701931 219085 701932
rect 222331 701996 222397 701997
rect 222331 701932 222332 701996
rect 222396 701932 222397 701996
rect 222331 701931 222397 701932
rect 219022 700501 219082 701931
rect 219019 700500 219085 700501
rect 219019 700436 219020 700500
rect 219084 700436 219085 700500
rect 219019 700435 219085 700436
rect 217712 687454 218032 687486
rect 217712 687218 217754 687454
rect 217990 687218 218032 687454
rect 217712 687134 218032 687218
rect 217712 686898 217754 687134
rect 217990 686898 218032 687134
rect 217712 686866 218032 686898
rect 217712 651454 218032 651486
rect 217712 651218 217754 651454
rect 217990 651218 218032 651454
rect 217712 651134 218032 651218
rect 217712 650898 217754 651134
rect 217990 650898 218032 651134
rect 217712 650866 218032 650898
rect 217712 615454 218032 615486
rect 217712 615218 217754 615454
rect 217990 615218 218032 615454
rect 217712 615134 218032 615218
rect 217712 614898 217754 615134
rect 217990 614898 218032 615134
rect 217712 614866 218032 614898
rect 217712 579454 218032 579486
rect 217712 579218 217754 579454
rect 217990 579218 218032 579454
rect 217712 579134 218032 579218
rect 217712 578898 217754 579134
rect 217990 578898 218032 579134
rect 217712 578866 218032 578898
rect 217712 543454 218032 543486
rect 217712 543218 217754 543454
rect 217990 543218 218032 543454
rect 217712 543134 218032 543218
rect 217712 542898 217754 543134
rect 217990 542898 218032 543134
rect 217712 542866 218032 542898
rect 217712 507454 218032 507486
rect 217712 507218 217754 507454
rect 217990 507218 218032 507454
rect 217712 507134 218032 507218
rect 217712 506898 217754 507134
rect 217990 506898 218032 507134
rect 217712 506866 218032 506898
rect 217712 471454 218032 471486
rect 217712 471218 217754 471454
rect 217990 471218 218032 471454
rect 217712 471134 218032 471218
rect 217712 470898 217754 471134
rect 217990 470898 218032 471134
rect 217712 470866 218032 470898
rect 217712 435454 218032 435486
rect 217712 435218 217754 435454
rect 217990 435218 218032 435454
rect 217712 435134 218032 435218
rect 217712 434898 217754 435134
rect 217990 434898 218032 435134
rect 217712 434866 218032 434898
rect 217712 399454 218032 399486
rect 217712 399218 217754 399454
rect 217990 399218 218032 399454
rect 217712 399134 218032 399218
rect 217712 398898 217754 399134
rect 217990 398898 218032 399134
rect 217712 398866 218032 398898
rect 217712 363454 218032 363486
rect 217712 363218 217754 363454
rect 217990 363218 218032 363454
rect 217712 363134 218032 363218
rect 217712 362898 217754 363134
rect 217990 362898 218032 363134
rect 217712 362866 218032 362898
rect 217712 327454 218032 327486
rect 217712 327218 217754 327454
rect 217990 327218 218032 327454
rect 217712 327134 218032 327218
rect 217712 326898 217754 327134
rect 217990 326898 218032 327134
rect 217712 326866 218032 326898
rect 217794 291454 218414 301784
rect 222334 300253 222394 701931
rect 222331 300252 222397 300253
rect 222331 300188 222332 300252
rect 222396 300188 222397 300252
rect 222331 300187 222397 300188
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 215339 125628 215405 125629
rect 215339 125564 215340 125628
rect 215404 125564 215405 125628
rect 215339 125563 215405 125564
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 212579 99516 212645 99517
rect 212579 99452 212580 99516
rect 212644 99452 212645 99516
rect 212579 99451 212645 99452
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 295174 222134 299784
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 298894 225854 299784
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 228774 244357 228834 702339
rect 229875 702268 229941 702269
rect 229875 702204 229876 702268
rect 229940 702204 229941 702268
rect 229875 702203 229941 702204
rect 229878 692790 229938 702203
rect 230059 701996 230125 701997
rect 230059 701932 230060 701996
rect 230124 701932 230125 701996
rect 230059 701931 230125 701932
rect 230243 701996 230309 701997
rect 230243 701932 230244 701996
rect 230308 701932 230309 701996
rect 230243 701931 230309 701932
rect 230062 699957 230122 701931
rect 230059 699956 230125 699957
rect 230059 699892 230060 699956
rect 230124 699892 230125 699956
rect 230059 699891 230125 699892
rect 229878 692730 230122 692790
rect 230062 300117 230122 692730
rect 230059 300116 230125 300117
rect 230059 300052 230060 300116
rect 230124 300052 230125 300116
rect 230059 300051 230125 300052
rect 228954 266614 229574 299784
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228771 244356 228837 244357
rect 228771 244292 228772 244356
rect 228836 244292 228837 244356
rect 228771 244291 228837 244292
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 230246 205733 230306 701931
rect 235794 701784 236414 705242
rect 239514 703784 240134 707162
rect 243234 703784 243854 709082
rect 246954 703784 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 251219 702540 251285 702541
rect 251219 702476 251220 702540
rect 251284 702476 251285 702540
rect 251219 702475 251285 702476
rect 251222 700093 251282 702475
rect 253794 701784 254414 704282
rect 257514 703784 258134 706202
rect 261234 703784 261854 708122
rect 264954 703784 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 701784 272414 705242
rect 275514 703784 276134 707162
rect 279234 703784 279854 709082
rect 282954 703784 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 701784 290414 704282
rect 293514 703784 294134 706202
rect 297234 703784 297854 708122
rect 300954 703784 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 701784 308414 705242
rect 311514 703784 312134 707162
rect 315234 703784 315854 709082
rect 318954 703784 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 316171 703084 316237 703085
rect 316171 703020 316172 703084
rect 316236 703020 316237 703084
rect 316171 703019 316237 703020
rect 316174 702810 316234 703019
rect 315806 702750 316234 702810
rect 315806 700501 315866 702750
rect 316171 702540 316237 702541
rect 316171 702476 316172 702540
rect 316236 702476 316237 702540
rect 316171 702475 316237 702476
rect 316174 700501 316234 702475
rect 325794 701784 326414 704282
rect 329514 703784 330134 706202
rect 333234 703784 333854 708122
rect 336954 703784 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 329787 703356 329853 703357
rect 329787 703292 329788 703356
rect 329852 703292 329853 703356
rect 329787 703291 329853 703292
rect 329790 701450 329850 703291
rect 343587 703220 343653 703221
rect 343587 703156 343588 703220
rect 343652 703156 343653 703220
rect 343587 703155 343653 703156
rect 333283 702540 333349 702541
rect 333283 702476 333284 702540
rect 333348 702476 333349 702540
rect 333283 702475 333349 702476
rect 329606 701390 329850 701450
rect 329606 701045 329666 701390
rect 333286 701045 333346 702475
rect 329603 701044 329669 701045
rect 329603 700980 329604 701044
rect 329668 700980 329669 701044
rect 329603 700979 329669 700980
rect 333283 701044 333349 701045
rect 333283 700980 333284 701044
rect 333348 700980 333349 701044
rect 333283 700979 333349 700980
rect 343590 700773 343650 703155
rect 343794 701784 344414 705242
rect 347514 703784 348134 707162
rect 351234 703784 351854 709082
rect 354954 703784 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 347819 703492 347885 703493
rect 347819 703428 347820 703492
rect 347884 703428 347885 703492
rect 347819 703427 347885 703428
rect 361435 703492 361501 703493
rect 361435 703428 361436 703492
rect 361500 703428 361501 703492
rect 361435 703427 361501 703428
rect 347822 702541 347882 703427
rect 345979 702540 346045 702541
rect 345979 702476 345980 702540
rect 346044 702476 346045 702540
rect 345979 702475 346045 702476
rect 347819 702540 347885 702541
rect 347819 702476 347820 702540
rect 347884 702476 347885 702540
rect 347819 702475 347885 702476
rect 352971 702540 353037 702541
rect 352971 702476 352972 702540
rect 353036 702476 353037 702540
rect 352971 702475 353037 702476
rect 345982 700773 346042 702475
rect 343587 700772 343653 700773
rect 343587 700708 343588 700772
rect 343652 700708 343653 700772
rect 343587 700707 343653 700708
rect 345979 700772 346045 700773
rect 345979 700708 345980 700772
rect 346044 700708 346045 700772
rect 345979 700707 346045 700708
rect 315803 700500 315869 700501
rect 315803 700436 315804 700500
rect 315868 700436 315869 700500
rect 315803 700435 315869 700436
rect 316171 700500 316237 700501
rect 316171 700436 316172 700500
rect 316236 700436 316237 700500
rect 316171 700435 316237 700436
rect 251219 700092 251285 700093
rect 251219 700028 251220 700092
rect 251284 700028 251285 700092
rect 251219 700027 251285 700028
rect 352974 699685 353034 702475
rect 361438 700637 361498 703427
rect 361794 701784 362414 704282
rect 365514 703784 366134 706202
rect 369234 703784 369854 708122
rect 372954 703784 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 365667 703084 365733 703085
rect 365667 703020 365668 703084
rect 365732 703020 365733 703084
rect 365667 703019 365733 703020
rect 365670 700773 365730 703019
rect 374867 702812 374933 702813
rect 374867 702748 374868 702812
rect 374932 702748 374933 702812
rect 374867 702747 374933 702748
rect 375419 702812 375485 702813
rect 375419 702748 375420 702812
rect 375484 702748 375485 702812
rect 375419 702747 375485 702748
rect 365851 702540 365917 702541
rect 365851 702476 365852 702540
rect 365916 702476 365917 702540
rect 365851 702475 365917 702476
rect 369715 702540 369781 702541
rect 369715 702476 369716 702540
rect 369780 702476 369781 702540
rect 369715 702475 369781 702476
rect 371923 702540 371989 702541
rect 371923 702476 371924 702540
rect 371988 702476 371989 702540
rect 371923 702475 371989 702476
rect 365667 700772 365733 700773
rect 365667 700708 365668 700772
rect 365732 700708 365733 700772
rect 365667 700707 365733 700708
rect 365854 700637 365914 702475
rect 369718 700773 369778 702475
rect 371926 701045 371986 702475
rect 374870 701045 374930 702747
rect 371923 701044 371989 701045
rect 371923 700980 371924 701044
rect 371988 700980 371989 701044
rect 371923 700979 371989 700980
rect 374867 701044 374933 701045
rect 374867 700980 374868 701044
rect 374932 700980 374933 701044
rect 374867 700979 374933 700980
rect 369715 700772 369781 700773
rect 369715 700708 369716 700772
rect 369780 700708 369781 700772
rect 369715 700707 369781 700708
rect 361435 700636 361501 700637
rect 361435 700572 361436 700636
rect 361500 700572 361501 700636
rect 361435 700571 361501 700572
rect 365851 700636 365917 700637
rect 365851 700572 365852 700636
rect 365916 700572 365917 700636
rect 365851 700571 365917 700572
rect 375422 699685 375482 702747
rect 378915 702540 378981 702541
rect 378915 702476 378916 702540
rect 378980 702476 378981 702540
rect 378915 702475 378981 702476
rect 378918 701045 378978 702475
rect 379794 701784 380414 705242
rect 383514 703784 384134 707162
rect 387234 703784 387854 709082
rect 390954 703784 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 391979 702676 392045 702677
rect 391979 702612 391980 702676
rect 392044 702612 392045 702676
rect 391979 702611 392045 702612
rect 391982 701045 392042 702611
rect 397794 701784 398414 704282
rect 401514 703784 402134 706202
rect 405234 703784 405854 708122
rect 408954 703784 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 412403 702676 412469 702677
rect 412403 702612 412404 702676
rect 412468 702612 412469 702676
rect 412403 702611 412469 702612
rect 378915 701044 378981 701045
rect 378915 700980 378916 701044
rect 378980 700980 378981 701044
rect 378915 700979 378981 700980
rect 391979 701044 392045 701045
rect 391979 700980 391980 701044
rect 392044 700980 392045 701044
rect 391979 700979 392045 700980
rect 412406 700909 412466 702611
rect 415794 701784 416414 705242
rect 419514 703784 420134 707162
rect 423234 703784 423854 709082
rect 426954 703784 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 427675 702676 427741 702677
rect 427675 702612 427676 702676
rect 427740 702612 427741 702676
rect 427675 702611 427741 702612
rect 427678 700909 427738 702611
rect 433794 701784 434414 704282
rect 437514 703784 438134 706202
rect 441234 703784 441854 708122
rect 444954 703784 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 701784 452414 705242
rect 455514 703784 456134 707162
rect 459234 703784 459854 709082
rect 462954 703784 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 701784 470414 704282
rect 473514 703784 474134 706202
rect 477234 703784 477854 708122
rect 480954 703784 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 701784 488414 705242
rect 491514 703784 492134 707162
rect 495234 703784 495854 709082
rect 498954 703784 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 701784 506414 704282
rect 509514 703784 510134 706202
rect 513234 703784 513854 708122
rect 516954 703784 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 701784 524414 705242
rect 527514 703784 528134 707162
rect 531234 703784 531854 709082
rect 534954 703784 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 701784 542414 704282
rect 545514 703784 546134 706202
rect 549234 703784 549854 708122
rect 552954 703784 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 701784 560414 705242
rect 563514 703784 564134 707162
rect 567234 703784 567854 709082
rect 570954 703784 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577451 703628 577517 703629
rect 577451 703564 577452 703628
rect 577516 703564 577517 703628
rect 577451 703563 577517 703564
rect 577267 703492 577333 703493
rect 577267 703428 577268 703492
rect 577332 703428 577333 703492
rect 577267 703427 577333 703428
rect 503483 701588 503549 701589
rect 503483 701524 503484 701588
rect 503548 701524 503549 701588
rect 503483 701523 503549 701524
rect 412403 700908 412469 700909
rect 412403 700844 412404 700908
rect 412468 700844 412469 700908
rect 412403 700843 412469 700844
rect 427675 700908 427741 700909
rect 427675 700844 427676 700908
rect 427740 700844 427741 700908
rect 427675 700843 427741 700844
rect 503486 700229 503546 701523
rect 510659 701180 510725 701181
rect 510659 701116 510660 701180
rect 510724 701116 510725 701180
rect 510659 701115 510725 701116
rect 520227 701180 520293 701181
rect 520227 701116 520228 701180
rect 520292 701116 520293 701180
rect 520227 701115 520293 701116
rect 528139 701180 528205 701181
rect 528139 701116 528140 701180
rect 528204 701116 528205 701180
rect 528139 701115 528205 701116
rect 532003 701180 532069 701181
rect 532003 701116 532004 701180
rect 532068 701116 532069 701180
rect 532003 701115 532069 701116
rect 532187 701180 532253 701181
rect 532187 701116 532188 701180
rect 532252 701116 532253 701180
rect 532187 701115 532253 701116
rect 545067 701180 545133 701181
rect 545067 701116 545068 701180
rect 545132 701116 545133 701180
rect 545067 701115 545133 701116
rect 550035 701180 550101 701181
rect 550035 701116 550036 701180
rect 550100 701116 550101 701180
rect 550035 701115 550101 701116
rect 559787 701180 559853 701181
rect 559787 701116 559788 701180
rect 559852 701116 559853 701180
rect 559787 701115 559853 701116
rect 570091 701180 570157 701181
rect 570091 701116 570092 701180
rect 570156 701116 570157 701180
rect 570091 701115 570157 701116
rect 572667 701180 572733 701181
rect 572667 701116 572668 701180
rect 572732 701116 572733 701180
rect 572667 701115 572733 701116
rect 503483 700228 503549 700229
rect 503483 700164 503484 700228
rect 503548 700164 503549 700228
rect 503483 700163 503549 700164
rect 352971 699684 353037 699685
rect 352971 699620 352972 699684
rect 353036 699620 353037 699684
rect 352971 699619 353037 699620
rect 375419 699684 375485 699685
rect 375419 699620 375420 699684
rect 375484 699620 375485 699684
rect 375419 699619 375485 699620
rect 248432 687454 248752 687486
rect 248432 687218 248474 687454
rect 248710 687218 248752 687454
rect 248432 687134 248752 687218
rect 248432 686898 248474 687134
rect 248710 686898 248752 687134
rect 248432 686866 248752 686898
rect 279152 687454 279472 687486
rect 279152 687218 279194 687454
rect 279430 687218 279472 687454
rect 279152 687134 279472 687218
rect 279152 686898 279194 687134
rect 279430 686898 279472 687134
rect 279152 686866 279472 686898
rect 309872 687454 310192 687486
rect 309872 687218 309914 687454
rect 310150 687218 310192 687454
rect 309872 687134 310192 687218
rect 309872 686898 309914 687134
rect 310150 686898 310192 687134
rect 309872 686866 310192 686898
rect 340592 687454 340912 687486
rect 340592 687218 340634 687454
rect 340870 687218 340912 687454
rect 340592 687134 340912 687218
rect 340592 686898 340634 687134
rect 340870 686898 340912 687134
rect 340592 686866 340912 686898
rect 371312 687454 371632 687486
rect 371312 687218 371354 687454
rect 371590 687218 371632 687454
rect 371312 687134 371632 687218
rect 371312 686898 371354 687134
rect 371590 686898 371632 687134
rect 371312 686866 371632 686898
rect 402032 687454 402352 687486
rect 402032 687218 402074 687454
rect 402310 687218 402352 687454
rect 402032 687134 402352 687218
rect 402032 686898 402074 687134
rect 402310 686898 402352 687134
rect 402032 686866 402352 686898
rect 432752 687454 433072 687486
rect 432752 687218 432794 687454
rect 433030 687218 433072 687454
rect 432752 687134 433072 687218
rect 432752 686898 432794 687134
rect 433030 686898 433072 687134
rect 432752 686866 433072 686898
rect 463472 687454 463792 687486
rect 463472 687218 463514 687454
rect 463750 687218 463792 687454
rect 463472 687134 463792 687218
rect 463472 686898 463514 687134
rect 463750 686898 463792 687134
rect 463472 686866 463792 686898
rect 494192 687454 494512 687486
rect 494192 687218 494234 687454
rect 494470 687218 494512 687454
rect 494192 687134 494512 687218
rect 494192 686898 494234 687134
rect 494470 686898 494512 687134
rect 494192 686866 494512 686898
rect 233072 669454 233392 669486
rect 233072 669218 233114 669454
rect 233350 669218 233392 669454
rect 233072 669134 233392 669218
rect 233072 668898 233114 669134
rect 233350 668898 233392 669134
rect 233072 668866 233392 668898
rect 263792 669454 264112 669486
rect 263792 669218 263834 669454
rect 264070 669218 264112 669454
rect 263792 669134 264112 669218
rect 263792 668898 263834 669134
rect 264070 668898 264112 669134
rect 263792 668866 264112 668898
rect 294512 669454 294832 669486
rect 294512 669218 294554 669454
rect 294790 669218 294832 669454
rect 294512 669134 294832 669218
rect 294512 668898 294554 669134
rect 294790 668898 294832 669134
rect 294512 668866 294832 668898
rect 325232 669454 325552 669486
rect 325232 669218 325274 669454
rect 325510 669218 325552 669454
rect 325232 669134 325552 669218
rect 325232 668898 325274 669134
rect 325510 668898 325552 669134
rect 325232 668866 325552 668898
rect 355952 669454 356272 669486
rect 355952 669218 355994 669454
rect 356230 669218 356272 669454
rect 355952 669134 356272 669218
rect 355952 668898 355994 669134
rect 356230 668898 356272 669134
rect 355952 668866 356272 668898
rect 386672 669454 386992 669486
rect 386672 669218 386714 669454
rect 386950 669218 386992 669454
rect 386672 669134 386992 669218
rect 386672 668898 386714 669134
rect 386950 668898 386992 669134
rect 386672 668866 386992 668898
rect 417392 669454 417712 669486
rect 417392 669218 417434 669454
rect 417670 669218 417712 669454
rect 417392 669134 417712 669218
rect 417392 668898 417434 669134
rect 417670 668898 417712 669134
rect 417392 668866 417712 668898
rect 448112 669454 448432 669486
rect 448112 669218 448154 669454
rect 448390 669218 448432 669454
rect 448112 669134 448432 669218
rect 448112 668898 448154 669134
rect 448390 668898 448432 669134
rect 448112 668866 448432 668898
rect 478832 669454 479152 669486
rect 478832 669218 478874 669454
rect 479110 669218 479152 669454
rect 478832 669134 479152 669218
rect 478832 668898 478874 669134
rect 479110 668898 479152 669134
rect 478832 668866 479152 668898
rect 509552 669454 509872 669486
rect 509552 669218 509594 669454
rect 509830 669218 509872 669454
rect 509552 669134 509872 669218
rect 509552 668898 509594 669134
rect 509830 668898 509872 669134
rect 509552 668866 509872 668898
rect 248432 651454 248752 651486
rect 248432 651218 248474 651454
rect 248710 651218 248752 651454
rect 248432 651134 248752 651218
rect 248432 650898 248474 651134
rect 248710 650898 248752 651134
rect 248432 650866 248752 650898
rect 279152 651454 279472 651486
rect 279152 651218 279194 651454
rect 279430 651218 279472 651454
rect 279152 651134 279472 651218
rect 279152 650898 279194 651134
rect 279430 650898 279472 651134
rect 279152 650866 279472 650898
rect 309872 651454 310192 651486
rect 309872 651218 309914 651454
rect 310150 651218 310192 651454
rect 309872 651134 310192 651218
rect 309872 650898 309914 651134
rect 310150 650898 310192 651134
rect 309872 650866 310192 650898
rect 340592 651454 340912 651486
rect 340592 651218 340634 651454
rect 340870 651218 340912 651454
rect 340592 651134 340912 651218
rect 340592 650898 340634 651134
rect 340870 650898 340912 651134
rect 340592 650866 340912 650898
rect 371312 651454 371632 651486
rect 371312 651218 371354 651454
rect 371590 651218 371632 651454
rect 371312 651134 371632 651218
rect 371312 650898 371354 651134
rect 371590 650898 371632 651134
rect 371312 650866 371632 650898
rect 402032 651454 402352 651486
rect 402032 651218 402074 651454
rect 402310 651218 402352 651454
rect 402032 651134 402352 651218
rect 402032 650898 402074 651134
rect 402310 650898 402352 651134
rect 402032 650866 402352 650898
rect 432752 651454 433072 651486
rect 432752 651218 432794 651454
rect 433030 651218 433072 651454
rect 432752 651134 433072 651218
rect 432752 650898 432794 651134
rect 433030 650898 433072 651134
rect 432752 650866 433072 650898
rect 463472 651454 463792 651486
rect 463472 651218 463514 651454
rect 463750 651218 463792 651454
rect 463472 651134 463792 651218
rect 463472 650898 463514 651134
rect 463750 650898 463792 651134
rect 463472 650866 463792 650898
rect 494192 651454 494512 651486
rect 494192 651218 494234 651454
rect 494470 651218 494512 651454
rect 494192 651134 494512 651218
rect 494192 650898 494234 651134
rect 494470 650898 494512 651134
rect 494192 650866 494512 650898
rect 233072 633454 233392 633486
rect 233072 633218 233114 633454
rect 233350 633218 233392 633454
rect 233072 633134 233392 633218
rect 233072 632898 233114 633134
rect 233350 632898 233392 633134
rect 233072 632866 233392 632898
rect 263792 633454 264112 633486
rect 263792 633218 263834 633454
rect 264070 633218 264112 633454
rect 263792 633134 264112 633218
rect 263792 632898 263834 633134
rect 264070 632898 264112 633134
rect 263792 632866 264112 632898
rect 294512 633454 294832 633486
rect 294512 633218 294554 633454
rect 294790 633218 294832 633454
rect 294512 633134 294832 633218
rect 294512 632898 294554 633134
rect 294790 632898 294832 633134
rect 294512 632866 294832 632898
rect 325232 633454 325552 633486
rect 325232 633218 325274 633454
rect 325510 633218 325552 633454
rect 325232 633134 325552 633218
rect 325232 632898 325274 633134
rect 325510 632898 325552 633134
rect 325232 632866 325552 632898
rect 355952 633454 356272 633486
rect 355952 633218 355994 633454
rect 356230 633218 356272 633454
rect 355952 633134 356272 633218
rect 355952 632898 355994 633134
rect 356230 632898 356272 633134
rect 355952 632866 356272 632898
rect 386672 633454 386992 633486
rect 386672 633218 386714 633454
rect 386950 633218 386992 633454
rect 386672 633134 386992 633218
rect 386672 632898 386714 633134
rect 386950 632898 386992 633134
rect 386672 632866 386992 632898
rect 417392 633454 417712 633486
rect 417392 633218 417434 633454
rect 417670 633218 417712 633454
rect 417392 633134 417712 633218
rect 417392 632898 417434 633134
rect 417670 632898 417712 633134
rect 417392 632866 417712 632898
rect 448112 633454 448432 633486
rect 448112 633218 448154 633454
rect 448390 633218 448432 633454
rect 448112 633134 448432 633218
rect 448112 632898 448154 633134
rect 448390 632898 448432 633134
rect 448112 632866 448432 632898
rect 478832 633454 479152 633486
rect 478832 633218 478874 633454
rect 479110 633218 479152 633454
rect 478832 633134 479152 633218
rect 478832 632898 478874 633134
rect 479110 632898 479152 633134
rect 478832 632866 479152 632898
rect 509552 633454 509872 633486
rect 509552 633218 509594 633454
rect 509830 633218 509872 633454
rect 509552 633134 509872 633218
rect 509552 632898 509594 633134
rect 509830 632898 509872 633134
rect 509552 632866 509872 632898
rect 248432 615454 248752 615486
rect 248432 615218 248474 615454
rect 248710 615218 248752 615454
rect 248432 615134 248752 615218
rect 248432 614898 248474 615134
rect 248710 614898 248752 615134
rect 248432 614866 248752 614898
rect 279152 615454 279472 615486
rect 279152 615218 279194 615454
rect 279430 615218 279472 615454
rect 279152 615134 279472 615218
rect 279152 614898 279194 615134
rect 279430 614898 279472 615134
rect 279152 614866 279472 614898
rect 309872 615454 310192 615486
rect 309872 615218 309914 615454
rect 310150 615218 310192 615454
rect 309872 615134 310192 615218
rect 309872 614898 309914 615134
rect 310150 614898 310192 615134
rect 309872 614866 310192 614898
rect 340592 615454 340912 615486
rect 340592 615218 340634 615454
rect 340870 615218 340912 615454
rect 340592 615134 340912 615218
rect 340592 614898 340634 615134
rect 340870 614898 340912 615134
rect 340592 614866 340912 614898
rect 371312 615454 371632 615486
rect 371312 615218 371354 615454
rect 371590 615218 371632 615454
rect 371312 615134 371632 615218
rect 371312 614898 371354 615134
rect 371590 614898 371632 615134
rect 371312 614866 371632 614898
rect 402032 615454 402352 615486
rect 402032 615218 402074 615454
rect 402310 615218 402352 615454
rect 402032 615134 402352 615218
rect 402032 614898 402074 615134
rect 402310 614898 402352 615134
rect 402032 614866 402352 614898
rect 432752 615454 433072 615486
rect 432752 615218 432794 615454
rect 433030 615218 433072 615454
rect 432752 615134 433072 615218
rect 432752 614898 432794 615134
rect 433030 614898 433072 615134
rect 432752 614866 433072 614898
rect 463472 615454 463792 615486
rect 463472 615218 463514 615454
rect 463750 615218 463792 615454
rect 463472 615134 463792 615218
rect 463472 614898 463514 615134
rect 463750 614898 463792 615134
rect 463472 614866 463792 614898
rect 494192 615454 494512 615486
rect 494192 615218 494234 615454
rect 494470 615218 494512 615454
rect 494192 615134 494512 615218
rect 494192 614898 494234 615134
rect 494470 614898 494512 615134
rect 494192 614866 494512 614898
rect 233072 597454 233392 597486
rect 233072 597218 233114 597454
rect 233350 597218 233392 597454
rect 233072 597134 233392 597218
rect 233072 596898 233114 597134
rect 233350 596898 233392 597134
rect 233072 596866 233392 596898
rect 263792 597454 264112 597486
rect 263792 597218 263834 597454
rect 264070 597218 264112 597454
rect 263792 597134 264112 597218
rect 263792 596898 263834 597134
rect 264070 596898 264112 597134
rect 263792 596866 264112 596898
rect 294512 597454 294832 597486
rect 294512 597218 294554 597454
rect 294790 597218 294832 597454
rect 294512 597134 294832 597218
rect 294512 596898 294554 597134
rect 294790 596898 294832 597134
rect 294512 596866 294832 596898
rect 325232 597454 325552 597486
rect 325232 597218 325274 597454
rect 325510 597218 325552 597454
rect 325232 597134 325552 597218
rect 325232 596898 325274 597134
rect 325510 596898 325552 597134
rect 325232 596866 325552 596898
rect 355952 597454 356272 597486
rect 355952 597218 355994 597454
rect 356230 597218 356272 597454
rect 355952 597134 356272 597218
rect 355952 596898 355994 597134
rect 356230 596898 356272 597134
rect 355952 596866 356272 596898
rect 386672 597454 386992 597486
rect 386672 597218 386714 597454
rect 386950 597218 386992 597454
rect 386672 597134 386992 597218
rect 386672 596898 386714 597134
rect 386950 596898 386992 597134
rect 386672 596866 386992 596898
rect 417392 597454 417712 597486
rect 417392 597218 417434 597454
rect 417670 597218 417712 597454
rect 417392 597134 417712 597218
rect 417392 596898 417434 597134
rect 417670 596898 417712 597134
rect 417392 596866 417712 596898
rect 448112 597454 448432 597486
rect 448112 597218 448154 597454
rect 448390 597218 448432 597454
rect 448112 597134 448432 597218
rect 448112 596898 448154 597134
rect 448390 596898 448432 597134
rect 448112 596866 448432 596898
rect 478832 597454 479152 597486
rect 478832 597218 478874 597454
rect 479110 597218 479152 597454
rect 478832 597134 479152 597218
rect 478832 596898 478874 597134
rect 479110 596898 479152 597134
rect 478832 596866 479152 596898
rect 509552 597454 509872 597486
rect 509552 597218 509594 597454
rect 509830 597218 509872 597454
rect 509552 597134 509872 597218
rect 509552 596898 509594 597134
rect 509830 596898 509872 597134
rect 509552 596866 509872 596898
rect 248432 579454 248752 579486
rect 248432 579218 248474 579454
rect 248710 579218 248752 579454
rect 248432 579134 248752 579218
rect 248432 578898 248474 579134
rect 248710 578898 248752 579134
rect 248432 578866 248752 578898
rect 279152 579454 279472 579486
rect 279152 579218 279194 579454
rect 279430 579218 279472 579454
rect 279152 579134 279472 579218
rect 279152 578898 279194 579134
rect 279430 578898 279472 579134
rect 279152 578866 279472 578898
rect 309872 579454 310192 579486
rect 309872 579218 309914 579454
rect 310150 579218 310192 579454
rect 309872 579134 310192 579218
rect 309872 578898 309914 579134
rect 310150 578898 310192 579134
rect 309872 578866 310192 578898
rect 340592 579454 340912 579486
rect 340592 579218 340634 579454
rect 340870 579218 340912 579454
rect 340592 579134 340912 579218
rect 340592 578898 340634 579134
rect 340870 578898 340912 579134
rect 340592 578866 340912 578898
rect 371312 579454 371632 579486
rect 371312 579218 371354 579454
rect 371590 579218 371632 579454
rect 371312 579134 371632 579218
rect 371312 578898 371354 579134
rect 371590 578898 371632 579134
rect 371312 578866 371632 578898
rect 402032 579454 402352 579486
rect 402032 579218 402074 579454
rect 402310 579218 402352 579454
rect 402032 579134 402352 579218
rect 402032 578898 402074 579134
rect 402310 578898 402352 579134
rect 402032 578866 402352 578898
rect 432752 579454 433072 579486
rect 432752 579218 432794 579454
rect 433030 579218 433072 579454
rect 432752 579134 433072 579218
rect 432752 578898 432794 579134
rect 433030 578898 433072 579134
rect 432752 578866 433072 578898
rect 463472 579454 463792 579486
rect 463472 579218 463514 579454
rect 463750 579218 463792 579454
rect 463472 579134 463792 579218
rect 463472 578898 463514 579134
rect 463750 578898 463792 579134
rect 463472 578866 463792 578898
rect 494192 579454 494512 579486
rect 494192 579218 494234 579454
rect 494470 579218 494512 579454
rect 494192 579134 494512 579218
rect 494192 578898 494234 579134
rect 494470 578898 494512 579134
rect 494192 578866 494512 578898
rect 233072 561454 233392 561486
rect 233072 561218 233114 561454
rect 233350 561218 233392 561454
rect 233072 561134 233392 561218
rect 233072 560898 233114 561134
rect 233350 560898 233392 561134
rect 233072 560866 233392 560898
rect 263792 561454 264112 561486
rect 263792 561218 263834 561454
rect 264070 561218 264112 561454
rect 263792 561134 264112 561218
rect 263792 560898 263834 561134
rect 264070 560898 264112 561134
rect 263792 560866 264112 560898
rect 294512 561454 294832 561486
rect 294512 561218 294554 561454
rect 294790 561218 294832 561454
rect 294512 561134 294832 561218
rect 294512 560898 294554 561134
rect 294790 560898 294832 561134
rect 294512 560866 294832 560898
rect 325232 561454 325552 561486
rect 325232 561218 325274 561454
rect 325510 561218 325552 561454
rect 325232 561134 325552 561218
rect 325232 560898 325274 561134
rect 325510 560898 325552 561134
rect 325232 560866 325552 560898
rect 355952 561454 356272 561486
rect 355952 561218 355994 561454
rect 356230 561218 356272 561454
rect 355952 561134 356272 561218
rect 355952 560898 355994 561134
rect 356230 560898 356272 561134
rect 355952 560866 356272 560898
rect 386672 561454 386992 561486
rect 386672 561218 386714 561454
rect 386950 561218 386992 561454
rect 386672 561134 386992 561218
rect 386672 560898 386714 561134
rect 386950 560898 386992 561134
rect 386672 560866 386992 560898
rect 417392 561454 417712 561486
rect 417392 561218 417434 561454
rect 417670 561218 417712 561454
rect 417392 561134 417712 561218
rect 417392 560898 417434 561134
rect 417670 560898 417712 561134
rect 417392 560866 417712 560898
rect 448112 561454 448432 561486
rect 448112 561218 448154 561454
rect 448390 561218 448432 561454
rect 448112 561134 448432 561218
rect 448112 560898 448154 561134
rect 448390 560898 448432 561134
rect 448112 560866 448432 560898
rect 478832 561454 479152 561486
rect 478832 561218 478874 561454
rect 479110 561218 479152 561454
rect 478832 561134 479152 561218
rect 478832 560898 478874 561134
rect 479110 560898 479152 561134
rect 478832 560866 479152 560898
rect 509552 561454 509872 561486
rect 509552 561218 509594 561454
rect 509830 561218 509872 561454
rect 509552 561134 509872 561218
rect 509552 560898 509594 561134
rect 509830 560898 509872 561134
rect 509552 560866 509872 560898
rect 248432 543454 248752 543486
rect 248432 543218 248474 543454
rect 248710 543218 248752 543454
rect 248432 543134 248752 543218
rect 248432 542898 248474 543134
rect 248710 542898 248752 543134
rect 248432 542866 248752 542898
rect 279152 543454 279472 543486
rect 279152 543218 279194 543454
rect 279430 543218 279472 543454
rect 279152 543134 279472 543218
rect 279152 542898 279194 543134
rect 279430 542898 279472 543134
rect 279152 542866 279472 542898
rect 309872 543454 310192 543486
rect 309872 543218 309914 543454
rect 310150 543218 310192 543454
rect 309872 543134 310192 543218
rect 309872 542898 309914 543134
rect 310150 542898 310192 543134
rect 309872 542866 310192 542898
rect 340592 543454 340912 543486
rect 340592 543218 340634 543454
rect 340870 543218 340912 543454
rect 340592 543134 340912 543218
rect 340592 542898 340634 543134
rect 340870 542898 340912 543134
rect 340592 542866 340912 542898
rect 371312 543454 371632 543486
rect 371312 543218 371354 543454
rect 371590 543218 371632 543454
rect 371312 543134 371632 543218
rect 371312 542898 371354 543134
rect 371590 542898 371632 543134
rect 371312 542866 371632 542898
rect 402032 543454 402352 543486
rect 402032 543218 402074 543454
rect 402310 543218 402352 543454
rect 402032 543134 402352 543218
rect 402032 542898 402074 543134
rect 402310 542898 402352 543134
rect 402032 542866 402352 542898
rect 432752 543454 433072 543486
rect 432752 543218 432794 543454
rect 433030 543218 433072 543454
rect 432752 543134 433072 543218
rect 432752 542898 432794 543134
rect 433030 542898 433072 543134
rect 432752 542866 433072 542898
rect 463472 543454 463792 543486
rect 463472 543218 463514 543454
rect 463750 543218 463792 543454
rect 463472 543134 463792 543218
rect 463472 542898 463514 543134
rect 463750 542898 463792 543134
rect 463472 542866 463792 542898
rect 494192 543454 494512 543486
rect 494192 543218 494234 543454
rect 494470 543218 494512 543454
rect 494192 543134 494512 543218
rect 494192 542898 494234 543134
rect 494470 542898 494512 543134
rect 494192 542866 494512 542898
rect 233072 525454 233392 525486
rect 233072 525218 233114 525454
rect 233350 525218 233392 525454
rect 233072 525134 233392 525218
rect 233072 524898 233114 525134
rect 233350 524898 233392 525134
rect 233072 524866 233392 524898
rect 263792 525454 264112 525486
rect 263792 525218 263834 525454
rect 264070 525218 264112 525454
rect 263792 525134 264112 525218
rect 263792 524898 263834 525134
rect 264070 524898 264112 525134
rect 263792 524866 264112 524898
rect 294512 525454 294832 525486
rect 294512 525218 294554 525454
rect 294790 525218 294832 525454
rect 294512 525134 294832 525218
rect 294512 524898 294554 525134
rect 294790 524898 294832 525134
rect 294512 524866 294832 524898
rect 325232 525454 325552 525486
rect 325232 525218 325274 525454
rect 325510 525218 325552 525454
rect 325232 525134 325552 525218
rect 325232 524898 325274 525134
rect 325510 524898 325552 525134
rect 325232 524866 325552 524898
rect 355952 525454 356272 525486
rect 355952 525218 355994 525454
rect 356230 525218 356272 525454
rect 355952 525134 356272 525218
rect 355952 524898 355994 525134
rect 356230 524898 356272 525134
rect 355952 524866 356272 524898
rect 386672 525454 386992 525486
rect 386672 525218 386714 525454
rect 386950 525218 386992 525454
rect 386672 525134 386992 525218
rect 386672 524898 386714 525134
rect 386950 524898 386992 525134
rect 386672 524866 386992 524898
rect 417392 525454 417712 525486
rect 417392 525218 417434 525454
rect 417670 525218 417712 525454
rect 417392 525134 417712 525218
rect 417392 524898 417434 525134
rect 417670 524898 417712 525134
rect 417392 524866 417712 524898
rect 448112 525454 448432 525486
rect 448112 525218 448154 525454
rect 448390 525218 448432 525454
rect 448112 525134 448432 525218
rect 448112 524898 448154 525134
rect 448390 524898 448432 525134
rect 448112 524866 448432 524898
rect 478832 525454 479152 525486
rect 478832 525218 478874 525454
rect 479110 525218 479152 525454
rect 478832 525134 479152 525218
rect 478832 524898 478874 525134
rect 479110 524898 479152 525134
rect 478832 524866 479152 524898
rect 509552 525454 509872 525486
rect 509552 525218 509594 525454
rect 509830 525218 509872 525454
rect 509552 525134 509872 525218
rect 509552 524898 509594 525134
rect 509830 524898 509872 525134
rect 509552 524866 509872 524898
rect 248432 507454 248752 507486
rect 248432 507218 248474 507454
rect 248710 507218 248752 507454
rect 248432 507134 248752 507218
rect 248432 506898 248474 507134
rect 248710 506898 248752 507134
rect 248432 506866 248752 506898
rect 279152 507454 279472 507486
rect 279152 507218 279194 507454
rect 279430 507218 279472 507454
rect 279152 507134 279472 507218
rect 279152 506898 279194 507134
rect 279430 506898 279472 507134
rect 279152 506866 279472 506898
rect 309872 507454 310192 507486
rect 309872 507218 309914 507454
rect 310150 507218 310192 507454
rect 309872 507134 310192 507218
rect 309872 506898 309914 507134
rect 310150 506898 310192 507134
rect 309872 506866 310192 506898
rect 340592 507454 340912 507486
rect 340592 507218 340634 507454
rect 340870 507218 340912 507454
rect 340592 507134 340912 507218
rect 340592 506898 340634 507134
rect 340870 506898 340912 507134
rect 340592 506866 340912 506898
rect 371312 507454 371632 507486
rect 371312 507218 371354 507454
rect 371590 507218 371632 507454
rect 371312 507134 371632 507218
rect 371312 506898 371354 507134
rect 371590 506898 371632 507134
rect 371312 506866 371632 506898
rect 402032 507454 402352 507486
rect 402032 507218 402074 507454
rect 402310 507218 402352 507454
rect 402032 507134 402352 507218
rect 402032 506898 402074 507134
rect 402310 506898 402352 507134
rect 402032 506866 402352 506898
rect 432752 507454 433072 507486
rect 432752 507218 432794 507454
rect 433030 507218 433072 507454
rect 432752 507134 433072 507218
rect 432752 506898 432794 507134
rect 433030 506898 433072 507134
rect 432752 506866 433072 506898
rect 463472 507454 463792 507486
rect 463472 507218 463514 507454
rect 463750 507218 463792 507454
rect 463472 507134 463792 507218
rect 463472 506898 463514 507134
rect 463750 506898 463792 507134
rect 463472 506866 463792 506898
rect 494192 507454 494512 507486
rect 494192 507218 494234 507454
rect 494470 507218 494512 507454
rect 494192 507134 494512 507218
rect 494192 506898 494234 507134
rect 494470 506898 494512 507134
rect 494192 506866 494512 506898
rect 233072 489454 233392 489486
rect 233072 489218 233114 489454
rect 233350 489218 233392 489454
rect 233072 489134 233392 489218
rect 233072 488898 233114 489134
rect 233350 488898 233392 489134
rect 233072 488866 233392 488898
rect 263792 489454 264112 489486
rect 263792 489218 263834 489454
rect 264070 489218 264112 489454
rect 263792 489134 264112 489218
rect 263792 488898 263834 489134
rect 264070 488898 264112 489134
rect 263792 488866 264112 488898
rect 294512 489454 294832 489486
rect 294512 489218 294554 489454
rect 294790 489218 294832 489454
rect 294512 489134 294832 489218
rect 294512 488898 294554 489134
rect 294790 488898 294832 489134
rect 294512 488866 294832 488898
rect 325232 489454 325552 489486
rect 325232 489218 325274 489454
rect 325510 489218 325552 489454
rect 325232 489134 325552 489218
rect 325232 488898 325274 489134
rect 325510 488898 325552 489134
rect 325232 488866 325552 488898
rect 355952 489454 356272 489486
rect 355952 489218 355994 489454
rect 356230 489218 356272 489454
rect 355952 489134 356272 489218
rect 355952 488898 355994 489134
rect 356230 488898 356272 489134
rect 355952 488866 356272 488898
rect 386672 489454 386992 489486
rect 386672 489218 386714 489454
rect 386950 489218 386992 489454
rect 386672 489134 386992 489218
rect 386672 488898 386714 489134
rect 386950 488898 386992 489134
rect 386672 488866 386992 488898
rect 417392 489454 417712 489486
rect 417392 489218 417434 489454
rect 417670 489218 417712 489454
rect 417392 489134 417712 489218
rect 417392 488898 417434 489134
rect 417670 488898 417712 489134
rect 417392 488866 417712 488898
rect 448112 489454 448432 489486
rect 448112 489218 448154 489454
rect 448390 489218 448432 489454
rect 448112 489134 448432 489218
rect 448112 488898 448154 489134
rect 448390 488898 448432 489134
rect 448112 488866 448432 488898
rect 478832 489454 479152 489486
rect 478832 489218 478874 489454
rect 479110 489218 479152 489454
rect 478832 489134 479152 489218
rect 478832 488898 478874 489134
rect 479110 488898 479152 489134
rect 478832 488866 479152 488898
rect 509552 489454 509872 489486
rect 509552 489218 509594 489454
rect 509830 489218 509872 489454
rect 509552 489134 509872 489218
rect 509552 488898 509594 489134
rect 509830 488898 509872 489134
rect 509552 488866 509872 488898
rect 248432 471454 248752 471486
rect 248432 471218 248474 471454
rect 248710 471218 248752 471454
rect 248432 471134 248752 471218
rect 248432 470898 248474 471134
rect 248710 470898 248752 471134
rect 248432 470866 248752 470898
rect 279152 471454 279472 471486
rect 279152 471218 279194 471454
rect 279430 471218 279472 471454
rect 279152 471134 279472 471218
rect 279152 470898 279194 471134
rect 279430 470898 279472 471134
rect 279152 470866 279472 470898
rect 309872 471454 310192 471486
rect 309872 471218 309914 471454
rect 310150 471218 310192 471454
rect 309872 471134 310192 471218
rect 309872 470898 309914 471134
rect 310150 470898 310192 471134
rect 309872 470866 310192 470898
rect 340592 471454 340912 471486
rect 340592 471218 340634 471454
rect 340870 471218 340912 471454
rect 340592 471134 340912 471218
rect 340592 470898 340634 471134
rect 340870 470898 340912 471134
rect 340592 470866 340912 470898
rect 371312 471454 371632 471486
rect 371312 471218 371354 471454
rect 371590 471218 371632 471454
rect 371312 471134 371632 471218
rect 371312 470898 371354 471134
rect 371590 470898 371632 471134
rect 371312 470866 371632 470898
rect 402032 471454 402352 471486
rect 402032 471218 402074 471454
rect 402310 471218 402352 471454
rect 402032 471134 402352 471218
rect 402032 470898 402074 471134
rect 402310 470898 402352 471134
rect 402032 470866 402352 470898
rect 432752 471454 433072 471486
rect 432752 471218 432794 471454
rect 433030 471218 433072 471454
rect 432752 471134 433072 471218
rect 432752 470898 432794 471134
rect 433030 470898 433072 471134
rect 432752 470866 433072 470898
rect 463472 471454 463792 471486
rect 463472 471218 463514 471454
rect 463750 471218 463792 471454
rect 463472 471134 463792 471218
rect 463472 470898 463514 471134
rect 463750 470898 463792 471134
rect 463472 470866 463792 470898
rect 494192 471454 494512 471486
rect 494192 471218 494234 471454
rect 494470 471218 494512 471454
rect 494192 471134 494512 471218
rect 494192 470898 494234 471134
rect 494470 470898 494512 471134
rect 494192 470866 494512 470898
rect 233072 453454 233392 453486
rect 233072 453218 233114 453454
rect 233350 453218 233392 453454
rect 233072 453134 233392 453218
rect 233072 452898 233114 453134
rect 233350 452898 233392 453134
rect 233072 452866 233392 452898
rect 263792 453454 264112 453486
rect 263792 453218 263834 453454
rect 264070 453218 264112 453454
rect 263792 453134 264112 453218
rect 263792 452898 263834 453134
rect 264070 452898 264112 453134
rect 263792 452866 264112 452898
rect 294512 453454 294832 453486
rect 294512 453218 294554 453454
rect 294790 453218 294832 453454
rect 294512 453134 294832 453218
rect 294512 452898 294554 453134
rect 294790 452898 294832 453134
rect 294512 452866 294832 452898
rect 325232 453454 325552 453486
rect 325232 453218 325274 453454
rect 325510 453218 325552 453454
rect 325232 453134 325552 453218
rect 325232 452898 325274 453134
rect 325510 452898 325552 453134
rect 325232 452866 325552 452898
rect 355952 453454 356272 453486
rect 355952 453218 355994 453454
rect 356230 453218 356272 453454
rect 355952 453134 356272 453218
rect 355952 452898 355994 453134
rect 356230 452898 356272 453134
rect 355952 452866 356272 452898
rect 386672 453454 386992 453486
rect 386672 453218 386714 453454
rect 386950 453218 386992 453454
rect 386672 453134 386992 453218
rect 386672 452898 386714 453134
rect 386950 452898 386992 453134
rect 386672 452866 386992 452898
rect 417392 453454 417712 453486
rect 417392 453218 417434 453454
rect 417670 453218 417712 453454
rect 417392 453134 417712 453218
rect 417392 452898 417434 453134
rect 417670 452898 417712 453134
rect 417392 452866 417712 452898
rect 448112 453454 448432 453486
rect 448112 453218 448154 453454
rect 448390 453218 448432 453454
rect 448112 453134 448432 453218
rect 448112 452898 448154 453134
rect 448390 452898 448432 453134
rect 448112 452866 448432 452898
rect 478832 453454 479152 453486
rect 478832 453218 478874 453454
rect 479110 453218 479152 453454
rect 478832 453134 479152 453218
rect 478832 452898 478874 453134
rect 479110 452898 479152 453134
rect 478832 452866 479152 452898
rect 509552 453454 509872 453486
rect 509552 453218 509594 453454
rect 509830 453218 509872 453454
rect 509552 453134 509872 453218
rect 509552 452898 509594 453134
rect 509830 452898 509872 453134
rect 509552 452866 509872 452898
rect 248432 435454 248752 435486
rect 248432 435218 248474 435454
rect 248710 435218 248752 435454
rect 248432 435134 248752 435218
rect 248432 434898 248474 435134
rect 248710 434898 248752 435134
rect 248432 434866 248752 434898
rect 279152 435454 279472 435486
rect 279152 435218 279194 435454
rect 279430 435218 279472 435454
rect 279152 435134 279472 435218
rect 279152 434898 279194 435134
rect 279430 434898 279472 435134
rect 279152 434866 279472 434898
rect 309872 435454 310192 435486
rect 309872 435218 309914 435454
rect 310150 435218 310192 435454
rect 309872 435134 310192 435218
rect 309872 434898 309914 435134
rect 310150 434898 310192 435134
rect 309872 434866 310192 434898
rect 340592 435454 340912 435486
rect 340592 435218 340634 435454
rect 340870 435218 340912 435454
rect 340592 435134 340912 435218
rect 340592 434898 340634 435134
rect 340870 434898 340912 435134
rect 340592 434866 340912 434898
rect 371312 435454 371632 435486
rect 371312 435218 371354 435454
rect 371590 435218 371632 435454
rect 371312 435134 371632 435218
rect 371312 434898 371354 435134
rect 371590 434898 371632 435134
rect 371312 434866 371632 434898
rect 402032 435454 402352 435486
rect 402032 435218 402074 435454
rect 402310 435218 402352 435454
rect 402032 435134 402352 435218
rect 402032 434898 402074 435134
rect 402310 434898 402352 435134
rect 402032 434866 402352 434898
rect 432752 435454 433072 435486
rect 432752 435218 432794 435454
rect 433030 435218 433072 435454
rect 432752 435134 433072 435218
rect 432752 434898 432794 435134
rect 433030 434898 433072 435134
rect 432752 434866 433072 434898
rect 463472 435454 463792 435486
rect 463472 435218 463514 435454
rect 463750 435218 463792 435454
rect 463472 435134 463792 435218
rect 463472 434898 463514 435134
rect 463750 434898 463792 435134
rect 463472 434866 463792 434898
rect 494192 435454 494512 435486
rect 494192 435218 494234 435454
rect 494470 435218 494512 435454
rect 494192 435134 494512 435218
rect 494192 434898 494234 435134
rect 494470 434898 494512 435134
rect 494192 434866 494512 434898
rect 233072 417454 233392 417486
rect 233072 417218 233114 417454
rect 233350 417218 233392 417454
rect 233072 417134 233392 417218
rect 233072 416898 233114 417134
rect 233350 416898 233392 417134
rect 233072 416866 233392 416898
rect 263792 417454 264112 417486
rect 263792 417218 263834 417454
rect 264070 417218 264112 417454
rect 263792 417134 264112 417218
rect 263792 416898 263834 417134
rect 264070 416898 264112 417134
rect 263792 416866 264112 416898
rect 294512 417454 294832 417486
rect 294512 417218 294554 417454
rect 294790 417218 294832 417454
rect 294512 417134 294832 417218
rect 294512 416898 294554 417134
rect 294790 416898 294832 417134
rect 294512 416866 294832 416898
rect 325232 417454 325552 417486
rect 325232 417218 325274 417454
rect 325510 417218 325552 417454
rect 325232 417134 325552 417218
rect 325232 416898 325274 417134
rect 325510 416898 325552 417134
rect 325232 416866 325552 416898
rect 355952 417454 356272 417486
rect 355952 417218 355994 417454
rect 356230 417218 356272 417454
rect 355952 417134 356272 417218
rect 355952 416898 355994 417134
rect 356230 416898 356272 417134
rect 355952 416866 356272 416898
rect 386672 417454 386992 417486
rect 386672 417218 386714 417454
rect 386950 417218 386992 417454
rect 386672 417134 386992 417218
rect 386672 416898 386714 417134
rect 386950 416898 386992 417134
rect 386672 416866 386992 416898
rect 417392 417454 417712 417486
rect 417392 417218 417434 417454
rect 417670 417218 417712 417454
rect 417392 417134 417712 417218
rect 417392 416898 417434 417134
rect 417670 416898 417712 417134
rect 417392 416866 417712 416898
rect 448112 417454 448432 417486
rect 448112 417218 448154 417454
rect 448390 417218 448432 417454
rect 448112 417134 448432 417218
rect 448112 416898 448154 417134
rect 448390 416898 448432 417134
rect 448112 416866 448432 416898
rect 478832 417454 479152 417486
rect 478832 417218 478874 417454
rect 479110 417218 479152 417454
rect 478832 417134 479152 417218
rect 478832 416898 478874 417134
rect 479110 416898 479152 417134
rect 478832 416866 479152 416898
rect 509552 417454 509872 417486
rect 509552 417218 509594 417454
rect 509830 417218 509872 417454
rect 509552 417134 509872 417218
rect 509552 416898 509594 417134
rect 509830 416898 509872 417134
rect 509552 416866 509872 416898
rect 248432 399454 248752 399486
rect 248432 399218 248474 399454
rect 248710 399218 248752 399454
rect 248432 399134 248752 399218
rect 248432 398898 248474 399134
rect 248710 398898 248752 399134
rect 248432 398866 248752 398898
rect 279152 399454 279472 399486
rect 279152 399218 279194 399454
rect 279430 399218 279472 399454
rect 279152 399134 279472 399218
rect 279152 398898 279194 399134
rect 279430 398898 279472 399134
rect 279152 398866 279472 398898
rect 309872 399454 310192 399486
rect 309872 399218 309914 399454
rect 310150 399218 310192 399454
rect 309872 399134 310192 399218
rect 309872 398898 309914 399134
rect 310150 398898 310192 399134
rect 309872 398866 310192 398898
rect 340592 399454 340912 399486
rect 340592 399218 340634 399454
rect 340870 399218 340912 399454
rect 340592 399134 340912 399218
rect 340592 398898 340634 399134
rect 340870 398898 340912 399134
rect 340592 398866 340912 398898
rect 371312 399454 371632 399486
rect 371312 399218 371354 399454
rect 371590 399218 371632 399454
rect 371312 399134 371632 399218
rect 371312 398898 371354 399134
rect 371590 398898 371632 399134
rect 371312 398866 371632 398898
rect 402032 399454 402352 399486
rect 402032 399218 402074 399454
rect 402310 399218 402352 399454
rect 402032 399134 402352 399218
rect 402032 398898 402074 399134
rect 402310 398898 402352 399134
rect 402032 398866 402352 398898
rect 432752 399454 433072 399486
rect 432752 399218 432794 399454
rect 433030 399218 433072 399454
rect 432752 399134 433072 399218
rect 432752 398898 432794 399134
rect 433030 398898 433072 399134
rect 432752 398866 433072 398898
rect 463472 399454 463792 399486
rect 463472 399218 463514 399454
rect 463750 399218 463792 399454
rect 463472 399134 463792 399218
rect 463472 398898 463514 399134
rect 463750 398898 463792 399134
rect 463472 398866 463792 398898
rect 494192 399454 494512 399486
rect 494192 399218 494234 399454
rect 494470 399218 494512 399454
rect 494192 399134 494512 399218
rect 494192 398898 494234 399134
rect 494470 398898 494512 399134
rect 494192 398866 494512 398898
rect 233072 381454 233392 381486
rect 233072 381218 233114 381454
rect 233350 381218 233392 381454
rect 233072 381134 233392 381218
rect 233072 380898 233114 381134
rect 233350 380898 233392 381134
rect 233072 380866 233392 380898
rect 263792 381454 264112 381486
rect 263792 381218 263834 381454
rect 264070 381218 264112 381454
rect 263792 381134 264112 381218
rect 263792 380898 263834 381134
rect 264070 380898 264112 381134
rect 263792 380866 264112 380898
rect 294512 381454 294832 381486
rect 294512 381218 294554 381454
rect 294790 381218 294832 381454
rect 294512 381134 294832 381218
rect 294512 380898 294554 381134
rect 294790 380898 294832 381134
rect 294512 380866 294832 380898
rect 325232 381454 325552 381486
rect 325232 381218 325274 381454
rect 325510 381218 325552 381454
rect 325232 381134 325552 381218
rect 325232 380898 325274 381134
rect 325510 380898 325552 381134
rect 325232 380866 325552 380898
rect 355952 381454 356272 381486
rect 355952 381218 355994 381454
rect 356230 381218 356272 381454
rect 355952 381134 356272 381218
rect 355952 380898 355994 381134
rect 356230 380898 356272 381134
rect 355952 380866 356272 380898
rect 386672 381454 386992 381486
rect 386672 381218 386714 381454
rect 386950 381218 386992 381454
rect 386672 381134 386992 381218
rect 386672 380898 386714 381134
rect 386950 380898 386992 381134
rect 386672 380866 386992 380898
rect 417392 381454 417712 381486
rect 417392 381218 417434 381454
rect 417670 381218 417712 381454
rect 417392 381134 417712 381218
rect 417392 380898 417434 381134
rect 417670 380898 417712 381134
rect 417392 380866 417712 380898
rect 448112 381454 448432 381486
rect 448112 381218 448154 381454
rect 448390 381218 448432 381454
rect 448112 381134 448432 381218
rect 448112 380898 448154 381134
rect 448390 380898 448432 381134
rect 448112 380866 448432 380898
rect 478832 381454 479152 381486
rect 478832 381218 478874 381454
rect 479110 381218 479152 381454
rect 478832 381134 479152 381218
rect 478832 380898 478874 381134
rect 479110 380898 479152 381134
rect 478832 380866 479152 380898
rect 509552 381454 509872 381486
rect 509552 381218 509594 381454
rect 509830 381218 509872 381454
rect 509552 381134 509872 381218
rect 509552 380898 509594 381134
rect 509830 380898 509872 381134
rect 509552 380866 509872 380898
rect 248432 363454 248752 363486
rect 248432 363218 248474 363454
rect 248710 363218 248752 363454
rect 248432 363134 248752 363218
rect 248432 362898 248474 363134
rect 248710 362898 248752 363134
rect 248432 362866 248752 362898
rect 279152 363454 279472 363486
rect 279152 363218 279194 363454
rect 279430 363218 279472 363454
rect 279152 363134 279472 363218
rect 279152 362898 279194 363134
rect 279430 362898 279472 363134
rect 279152 362866 279472 362898
rect 309872 363454 310192 363486
rect 309872 363218 309914 363454
rect 310150 363218 310192 363454
rect 309872 363134 310192 363218
rect 309872 362898 309914 363134
rect 310150 362898 310192 363134
rect 309872 362866 310192 362898
rect 340592 363454 340912 363486
rect 340592 363218 340634 363454
rect 340870 363218 340912 363454
rect 340592 363134 340912 363218
rect 340592 362898 340634 363134
rect 340870 362898 340912 363134
rect 340592 362866 340912 362898
rect 371312 363454 371632 363486
rect 371312 363218 371354 363454
rect 371590 363218 371632 363454
rect 371312 363134 371632 363218
rect 371312 362898 371354 363134
rect 371590 362898 371632 363134
rect 371312 362866 371632 362898
rect 402032 363454 402352 363486
rect 402032 363218 402074 363454
rect 402310 363218 402352 363454
rect 402032 363134 402352 363218
rect 402032 362898 402074 363134
rect 402310 362898 402352 363134
rect 402032 362866 402352 362898
rect 432752 363454 433072 363486
rect 432752 363218 432794 363454
rect 433030 363218 433072 363454
rect 432752 363134 433072 363218
rect 432752 362898 432794 363134
rect 433030 362898 433072 363134
rect 432752 362866 433072 362898
rect 463472 363454 463792 363486
rect 463472 363218 463514 363454
rect 463750 363218 463792 363454
rect 463472 363134 463792 363218
rect 463472 362898 463514 363134
rect 463750 362898 463792 363134
rect 463472 362866 463792 362898
rect 494192 363454 494512 363486
rect 494192 363218 494234 363454
rect 494470 363218 494512 363454
rect 494192 363134 494512 363218
rect 494192 362898 494234 363134
rect 494470 362898 494512 363134
rect 494192 362866 494512 362898
rect 233072 345454 233392 345486
rect 233072 345218 233114 345454
rect 233350 345218 233392 345454
rect 233072 345134 233392 345218
rect 233072 344898 233114 345134
rect 233350 344898 233392 345134
rect 233072 344866 233392 344898
rect 263792 345454 264112 345486
rect 263792 345218 263834 345454
rect 264070 345218 264112 345454
rect 263792 345134 264112 345218
rect 263792 344898 263834 345134
rect 264070 344898 264112 345134
rect 263792 344866 264112 344898
rect 294512 345454 294832 345486
rect 294512 345218 294554 345454
rect 294790 345218 294832 345454
rect 294512 345134 294832 345218
rect 294512 344898 294554 345134
rect 294790 344898 294832 345134
rect 294512 344866 294832 344898
rect 325232 345454 325552 345486
rect 325232 345218 325274 345454
rect 325510 345218 325552 345454
rect 325232 345134 325552 345218
rect 325232 344898 325274 345134
rect 325510 344898 325552 345134
rect 325232 344866 325552 344898
rect 355952 345454 356272 345486
rect 355952 345218 355994 345454
rect 356230 345218 356272 345454
rect 355952 345134 356272 345218
rect 355952 344898 355994 345134
rect 356230 344898 356272 345134
rect 355952 344866 356272 344898
rect 386672 345454 386992 345486
rect 386672 345218 386714 345454
rect 386950 345218 386992 345454
rect 386672 345134 386992 345218
rect 386672 344898 386714 345134
rect 386950 344898 386992 345134
rect 386672 344866 386992 344898
rect 417392 345454 417712 345486
rect 417392 345218 417434 345454
rect 417670 345218 417712 345454
rect 417392 345134 417712 345218
rect 417392 344898 417434 345134
rect 417670 344898 417712 345134
rect 417392 344866 417712 344898
rect 448112 345454 448432 345486
rect 448112 345218 448154 345454
rect 448390 345218 448432 345454
rect 448112 345134 448432 345218
rect 448112 344898 448154 345134
rect 448390 344898 448432 345134
rect 448112 344866 448432 344898
rect 478832 345454 479152 345486
rect 478832 345218 478874 345454
rect 479110 345218 479152 345454
rect 478832 345134 479152 345218
rect 478832 344898 478874 345134
rect 479110 344898 479152 345134
rect 478832 344866 479152 344898
rect 509552 345454 509872 345486
rect 509552 345218 509594 345454
rect 509830 345218 509872 345454
rect 509552 345134 509872 345218
rect 509552 344898 509594 345134
rect 509830 344898 509872 345134
rect 509552 344866 509872 344898
rect 248432 327454 248752 327486
rect 248432 327218 248474 327454
rect 248710 327218 248752 327454
rect 248432 327134 248752 327218
rect 248432 326898 248474 327134
rect 248710 326898 248752 327134
rect 248432 326866 248752 326898
rect 279152 327454 279472 327486
rect 279152 327218 279194 327454
rect 279430 327218 279472 327454
rect 279152 327134 279472 327218
rect 279152 326898 279194 327134
rect 279430 326898 279472 327134
rect 279152 326866 279472 326898
rect 309872 327454 310192 327486
rect 309872 327218 309914 327454
rect 310150 327218 310192 327454
rect 309872 327134 310192 327218
rect 309872 326898 309914 327134
rect 310150 326898 310192 327134
rect 309872 326866 310192 326898
rect 340592 327454 340912 327486
rect 340592 327218 340634 327454
rect 340870 327218 340912 327454
rect 340592 327134 340912 327218
rect 340592 326898 340634 327134
rect 340870 326898 340912 327134
rect 340592 326866 340912 326898
rect 371312 327454 371632 327486
rect 371312 327218 371354 327454
rect 371590 327218 371632 327454
rect 371312 327134 371632 327218
rect 371312 326898 371354 327134
rect 371590 326898 371632 327134
rect 371312 326866 371632 326898
rect 402032 327454 402352 327486
rect 402032 327218 402074 327454
rect 402310 327218 402352 327454
rect 402032 327134 402352 327218
rect 402032 326898 402074 327134
rect 402310 326898 402352 327134
rect 402032 326866 402352 326898
rect 432752 327454 433072 327486
rect 432752 327218 432794 327454
rect 433030 327218 433072 327454
rect 432752 327134 433072 327218
rect 432752 326898 432794 327134
rect 433030 326898 433072 327134
rect 432752 326866 433072 326898
rect 463472 327454 463792 327486
rect 463472 327218 463514 327454
rect 463750 327218 463792 327454
rect 463472 327134 463792 327218
rect 463472 326898 463514 327134
rect 463750 326898 463792 327134
rect 463472 326866 463792 326898
rect 494192 327454 494512 327486
rect 494192 327218 494234 327454
rect 494470 327218 494512 327454
rect 494192 327134 494512 327218
rect 494192 326898 494234 327134
rect 494470 326898 494512 327134
rect 494192 326866 494512 326898
rect 233072 309454 233392 309486
rect 233072 309218 233114 309454
rect 233350 309218 233392 309454
rect 233072 309134 233392 309218
rect 233072 308898 233114 309134
rect 233350 308898 233392 309134
rect 233072 308866 233392 308898
rect 263792 309454 264112 309486
rect 263792 309218 263834 309454
rect 264070 309218 264112 309454
rect 263792 309134 264112 309218
rect 263792 308898 263834 309134
rect 264070 308898 264112 309134
rect 263792 308866 264112 308898
rect 294512 309454 294832 309486
rect 294512 309218 294554 309454
rect 294790 309218 294832 309454
rect 294512 309134 294832 309218
rect 294512 308898 294554 309134
rect 294790 308898 294832 309134
rect 294512 308866 294832 308898
rect 325232 309454 325552 309486
rect 325232 309218 325274 309454
rect 325510 309218 325552 309454
rect 325232 309134 325552 309218
rect 325232 308898 325274 309134
rect 325510 308898 325552 309134
rect 325232 308866 325552 308898
rect 355952 309454 356272 309486
rect 355952 309218 355994 309454
rect 356230 309218 356272 309454
rect 355952 309134 356272 309218
rect 355952 308898 355994 309134
rect 356230 308898 356272 309134
rect 355952 308866 356272 308898
rect 386672 309454 386992 309486
rect 386672 309218 386714 309454
rect 386950 309218 386992 309454
rect 386672 309134 386992 309218
rect 386672 308898 386714 309134
rect 386950 308898 386992 309134
rect 386672 308866 386992 308898
rect 417392 309454 417712 309486
rect 417392 309218 417434 309454
rect 417670 309218 417712 309454
rect 417392 309134 417712 309218
rect 417392 308898 417434 309134
rect 417670 308898 417712 309134
rect 417392 308866 417712 308898
rect 448112 309454 448432 309486
rect 448112 309218 448154 309454
rect 448390 309218 448432 309454
rect 448112 309134 448432 309218
rect 448112 308898 448154 309134
rect 448390 308898 448432 309134
rect 448112 308866 448432 308898
rect 478832 309454 479152 309486
rect 478832 309218 478874 309454
rect 479110 309218 479152 309454
rect 478832 309134 479152 309218
rect 478832 308898 478874 309134
rect 479110 308898 479152 309134
rect 478832 308866 479152 308898
rect 509552 309454 509872 309486
rect 509552 309218 509594 309454
rect 509830 309218 509872 309454
rect 509552 309134 509872 309218
rect 509552 308898 509594 309134
rect 509830 308898 509872 309134
rect 509552 308866 509872 308898
rect 510662 303517 510722 701115
rect 510659 303516 510725 303517
rect 510659 303452 510660 303516
rect 510724 303452 510725 303516
rect 510659 303451 510725 303452
rect 235794 273454 236414 301784
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 230243 205732 230309 205733
rect 230243 205668 230244 205732
rect 230308 205668 230309 205732
rect 230243 205667 230309 205668
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 277174 240134 299784
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 280894 243854 299784
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 284614 247574 299784
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 291454 254414 301784
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 295174 258134 299784
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 298894 261854 299784
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 266614 265574 299784
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 273454 272414 301784
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 277174 276134 299784
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 280894 279854 299784
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 284614 283574 299784
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 291454 290414 301784
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 295174 294134 299784
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 298894 297854 299784
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 266614 301574 299784
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 273454 308414 301784
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 277174 312134 299784
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 280894 315854 299784
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 284614 319574 299784
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 291454 326414 301784
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 295174 330134 299784
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 298894 333854 299784
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 266614 337574 299784
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 273454 344414 301784
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 277174 348134 299784
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 280894 351854 299784
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 284614 355574 299784
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 291454 362414 301784
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 295174 366134 299784
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 298894 369854 299784
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 266614 373574 299784
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 273454 380414 301784
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 277174 384134 299784
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 280894 387854 299784
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 284614 391574 299784
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 291454 398414 301784
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 295174 402134 299784
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 298894 405854 299784
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 266614 409574 299784
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 273454 416414 301784
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 277174 420134 299784
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 280894 423854 299784
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 284614 427574 299784
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 291454 434414 301784
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 295174 438134 299784
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 298894 441854 299784
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 266614 445574 299784
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 273454 452414 301784
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 277174 456134 299784
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 280894 459854 299784
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 284614 463574 299784
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 291454 470414 301784
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 295174 474134 299784
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 298894 477854 299784
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 266614 481574 299784
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 273454 488414 301784
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 277174 492134 299784
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 280894 495854 299784
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 284614 499574 299784
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 291454 506414 301784
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 295174 510134 299784
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 298894 513854 299784
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 266614 517574 299784
rect 520230 267749 520290 701115
rect 528142 699821 528202 701115
rect 528139 699820 528205 699821
rect 528139 699756 528140 699820
rect 528204 699756 528205 699820
rect 528139 699755 528205 699756
rect 524912 687454 525232 687486
rect 524912 687218 524954 687454
rect 525190 687218 525232 687454
rect 524912 687134 525232 687218
rect 524912 686898 524954 687134
rect 525190 686898 525232 687134
rect 524912 686866 525232 686898
rect 524912 651454 525232 651486
rect 524912 651218 524954 651454
rect 525190 651218 525232 651454
rect 524912 651134 525232 651218
rect 524912 650898 524954 651134
rect 525190 650898 525232 651134
rect 524912 650866 525232 650898
rect 524912 615454 525232 615486
rect 524912 615218 524954 615454
rect 525190 615218 525232 615454
rect 524912 615134 525232 615218
rect 524912 614898 524954 615134
rect 525190 614898 525232 615134
rect 524912 614866 525232 614898
rect 524912 579454 525232 579486
rect 524912 579218 524954 579454
rect 525190 579218 525232 579454
rect 524912 579134 525232 579218
rect 524912 578898 524954 579134
rect 525190 578898 525232 579134
rect 524912 578866 525232 578898
rect 524912 543454 525232 543486
rect 524912 543218 524954 543454
rect 525190 543218 525232 543454
rect 524912 543134 525232 543218
rect 524912 542898 524954 543134
rect 525190 542898 525232 543134
rect 524912 542866 525232 542898
rect 524912 507454 525232 507486
rect 524912 507218 524954 507454
rect 525190 507218 525232 507454
rect 524912 507134 525232 507218
rect 524912 506898 524954 507134
rect 525190 506898 525232 507134
rect 524912 506866 525232 506898
rect 524912 471454 525232 471486
rect 524912 471218 524954 471454
rect 525190 471218 525232 471454
rect 524912 471134 525232 471218
rect 524912 470898 524954 471134
rect 525190 470898 525232 471134
rect 524912 470866 525232 470898
rect 524912 435454 525232 435486
rect 524912 435218 524954 435454
rect 525190 435218 525232 435454
rect 524912 435134 525232 435218
rect 524912 434898 524954 435134
rect 525190 434898 525232 435134
rect 524912 434866 525232 434898
rect 524912 399454 525232 399486
rect 524912 399218 524954 399454
rect 525190 399218 525232 399454
rect 524912 399134 525232 399218
rect 524912 398898 524954 399134
rect 525190 398898 525232 399134
rect 524912 398866 525232 398898
rect 524912 363454 525232 363486
rect 524912 363218 524954 363454
rect 525190 363218 525232 363454
rect 524912 363134 525232 363218
rect 524912 362898 524954 363134
rect 525190 362898 525232 363134
rect 524912 362866 525232 362898
rect 524912 327454 525232 327486
rect 524912 327218 524954 327454
rect 525190 327218 525232 327454
rect 524912 327134 525232 327218
rect 524912 326898 524954 327134
rect 525190 326898 525232 327134
rect 524912 326866 525232 326898
rect 523794 273454 524414 301784
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 520227 267748 520293 267749
rect 520227 267684 520228 267748
rect 520292 267684 520293 267748
rect 520227 267683 520293 267684
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 277174 528134 299784
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 280894 531854 299784
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 532006 215253 532066 701115
rect 532190 700365 532250 701115
rect 532187 700364 532253 700365
rect 532187 700300 532188 700364
rect 532252 700300 532253 700364
rect 532187 700299 532253 700300
rect 540272 669454 540592 669486
rect 540272 669218 540314 669454
rect 540550 669218 540592 669454
rect 540272 669134 540592 669218
rect 540272 668898 540314 669134
rect 540550 668898 540592 669134
rect 540272 668866 540592 668898
rect 540272 633454 540592 633486
rect 540272 633218 540314 633454
rect 540550 633218 540592 633454
rect 540272 633134 540592 633218
rect 540272 632898 540314 633134
rect 540550 632898 540592 633134
rect 540272 632866 540592 632898
rect 540272 597454 540592 597486
rect 540272 597218 540314 597454
rect 540550 597218 540592 597454
rect 540272 597134 540592 597218
rect 540272 596898 540314 597134
rect 540550 596898 540592 597134
rect 540272 596866 540592 596898
rect 540272 561454 540592 561486
rect 540272 561218 540314 561454
rect 540550 561218 540592 561454
rect 540272 561134 540592 561218
rect 540272 560898 540314 561134
rect 540550 560898 540592 561134
rect 540272 560866 540592 560898
rect 540272 525454 540592 525486
rect 540272 525218 540314 525454
rect 540550 525218 540592 525454
rect 540272 525134 540592 525218
rect 540272 524898 540314 525134
rect 540550 524898 540592 525134
rect 540272 524866 540592 524898
rect 540272 489454 540592 489486
rect 540272 489218 540314 489454
rect 540550 489218 540592 489454
rect 540272 489134 540592 489218
rect 540272 488898 540314 489134
rect 540550 488898 540592 489134
rect 540272 488866 540592 488898
rect 540272 453454 540592 453486
rect 540272 453218 540314 453454
rect 540550 453218 540592 453454
rect 540272 453134 540592 453218
rect 540272 452898 540314 453134
rect 540550 452898 540592 453134
rect 540272 452866 540592 452898
rect 540272 417454 540592 417486
rect 540272 417218 540314 417454
rect 540550 417218 540592 417454
rect 540272 417134 540592 417218
rect 540272 416898 540314 417134
rect 540550 416898 540592 417134
rect 540272 416866 540592 416898
rect 540272 381454 540592 381486
rect 540272 381218 540314 381454
rect 540550 381218 540592 381454
rect 540272 381134 540592 381218
rect 540272 380898 540314 381134
rect 540550 380898 540592 381134
rect 540272 380866 540592 380898
rect 540272 345454 540592 345486
rect 540272 345218 540314 345454
rect 540550 345218 540592 345454
rect 540272 345134 540592 345218
rect 540272 344898 540314 345134
rect 540550 344898 540592 345134
rect 540272 344866 540592 344898
rect 540272 309454 540592 309486
rect 540272 309218 540314 309454
rect 540550 309218 540592 309454
rect 540272 309134 540592 309218
rect 540272 308898 540314 309134
rect 540550 308898 540592 309134
rect 540272 308866 540592 308898
rect 534954 284614 535574 299784
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 532003 215252 532069 215253
rect 532003 215188 532004 215252
rect 532068 215188 532069 215252
rect 532003 215187 532069 215188
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 291454 542414 301784
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 545070 138005 545130 701115
rect 545514 295174 546134 299784
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545067 138004 545133 138005
rect 545067 137940 545068 138004
rect 545132 137940 545133 138004
rect 545067 137939 545133 137940
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 298894 549854 299784
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 550038 150381 550098 701115
rect 559790 700501 559850 701115
rect 559787 700500 559853 700501
rect 559787 700436 559788 700500
rect 559852 700436 559853 700500
rect 559787 700435 559853 700436
rect 555632 687454 555952 687486
rect 555632 687218 555674 687454
rect 555910 687218 555952 687454
rect 555632 687134 555952 687218
rect 555632 686898 555674 687134
rect 555910 686898 555952 687134
rect 555632 686866 555952 686898
rect 555632 651454 555952 651486
rect 555632 651218 555674 651454
rect 555910 651218 555952 651454
rect 555632 651134 555952 651218
rect 555632 650898 555674 651134
rect 555910 650898 555952 651134
rect 555632 650866 555952 650898
rect 555632 615454 555952 615486
rect 555632 615218 555674 615454
rect 555910 615218 555952 615454
rect 555632 615134 555952 615218
rect 555632 614898 555674 615134
rect 555910 614898 555952 615134
rect 555632 614866 555952 614898
rect 555632 579454 555952 579486
rect 555632 579218 555674 579454
rect 555910 579218 555952 579454
rect 555632 579134 555952 579218
rect 555632 578898 555674 579134
rect 555910 578898 555952 579134
rect 555632 578866 555952 578898
rect 555632 543454 555952 543486
rect 555632 543218 555674 543454
rect 555910 543218 555952 543454
rect 555632 543134 555952 543218
rect 555632 542898 555674 543134
rect 555910 542898 555952 543134
rect 555632 542866 555952 542898
rect 555632 507454 555952 507486
rect 555632 507218 555674 507454
rect 555910 507218 555952 507454
rect 555632 507134 555952 507218
rect 555632 506898 555674 507134
rect 555910 506898 555952 507134
rect 555632 506866 555952 506898
rect 555632 471454 555952 471486
rect 555632 471218 555674 471454
rect 555910 471218 555952 471454
rect 555632 471134 555952 471218
rect 555632 470898 555674 471134
rect 555910 470898 555952 471134
rect 555632 470866 555952 470898
rect 555632 435454 555952 435486
rect 555632 435218 555674 435454
rect 555910 435218 555952 435454
rect 555632 435134 555952 435218
rect 555632 434898 555674 435134
rect 555910 434898 555952 435134
rect 555632 434866 555952 434898
rect 555632 399454 555952 399486
rect 555632 399218 555674 399454
rect 555910 399218 555952 399454
rect 555632 399134 555952 399218
rect 555632 398898 555674 399134
rect 555910 398898 555952 399134
rect 555632 398866 555952 398898
rect 555632 363454 555952 363486
rect 555632 363218 555674 363454
rect 555910 363218 555952 363454
rect 555632 363134 555952 363218
rect 555632 362898 555674 363134
rect 555910 362898 555952 363134
rect 555632 362866 555952 362898
rect 555632 327454 555952 327486
rect 555632 327218 555674 327454
rect 555910 327218 555952 327454
rect 555632 327134 555952 327218
rect 555632 326898 555674 327134
rect 555910 326898 555952 327134
rect 555632 326866 555952 326898
rect 552954 266614 553574 299784
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 550035 150380 550101 150381
rect 550035 150316 550036 150380
rect 550100 150316 550101 150380
rect 550035 150315 550101 150316
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 273454 560414 301784
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 277174 564134 299784
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 280894 567854 299784
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 570094 59261 570154 701115
rect 570992 669454 571312 669486
rect 570992 669218 571034 669454
rect 571270 669218 571312 669454
rect 570992 669134 571312 669218
rect 570992 668898 571034 669134
rect 571270 668898 571312 669134
rect 570992 668866 571312 668898
rect 570992 633454 571312 633486
rect 570992 633218 571034 633454
rect 571270 633218 571312 633454
rect 570992 633134 571312 633218
rect 570992 632898 571034 633134
rect 571270 632898 571312 633134
rect 570992 632866 571312 632898
rect 570992 597454 571312 597486
rect 570992 597218 571034 597454
rect 571270 597218 571312 597454
rect 570992 597134 571312 597218
rect 570992 596898 571034 597134
rect 571270 596898 571312 597134
rect 570992 596866 571312 596898
rect 570992 561454 571312 561486
rect 570992 561218 571034 561454
rect 571270 561218 571312 561454
rect 570992 561134 571312 561218
rect 570992 560898 571034 561134
rect 571270 560898 571312 561134
rect 570992 560866 571312 560898
rect 570992 525454 571312 525486
rect 570992 525218 571034 525454
rect 571270 525218 571312 525454
rect 570992 525134 571312 525218
rect 570992 524898 571034 525134
rect 571270 524898 571312 525134
rect 570992 524866 571312 524898
rect 570992 489454 571312 489486
rect 570992 489218 571034 489454
rect 571270 489218 571312 489454
rect 570992 489134 571312 489218
rect 570992 488898 571034 489134
rect 571270 488898 571312 489134
rect 570992 488866 571312 488898
rect 570992 453454 571312 453486
rect 570992 453218 571034 453454
rect 571270 453218 571312 453454
rect 570992 453134 571312 453218
rect 570992 452898 571034 453134
rect 571270 452898 571312 453134
rect 570992 452866 571312 452898
rect 570992 417454 571312 417486
rect 570992 417218 571034 417454
rect 571270 417218 571312 417454
rect 570992 417134 571312 417218
rect 570992 416898 571034 417134
rect 571270 416898 571312 417134
rect 570992 416866 571312 416898
rect 570992 381454 571312 381486
rect 570992 381218 571034 381454
rect 571270 381218 571312 381454
rect 570992 381134 571312 381218
rect 570992 380898 571034 381134
rect 571270 380898 571312 381134
rect 570992 380866 571312 380898
rect 570992 345454 571312 345486
rect 570992 345218 571034 345454
rect 571270 345218 571312 345454
rect 570992 345134 571312 345218
rect 570992 344898 571034 345134
rect 571270 344898 571312 345134
rect 570992 344866 571312 344898
rect 570992 309454 571312 309486
rect 570992 309218 571034 309454
rect 571270 309218 571312 309454
rect 570992 309134 571312 309218
rect 570992 308898 571034 309134
rect 571270 308898 571312 309134
rect 570992 308866 571312 308898
rect 570954 284614 571574 299784
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570091 59260 570157 59261
rect 570091 59196 570092 59260
rect 570156 59196 570157 59260
rect 570091 59195 570157 59196
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 32614 571574 68058
rect 572670 33149 572730 701115
rect 577270 364350 577330 703427
rect 577454 576870 577514 703563
rect 577635 703084 577701 703085
rect 577635 703020 577636 703084
rect 577700 703020 577701 703084
rect 577635 703019 577701 703020
rect 577638 634830 577698 703019
rect 577794 701784 578414 704282
rect 581514 703784 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 580579 703220 580645 703221
rect 580579 703156 580580 703220
rect 580644 703156 580645 703220
rect 580579 703155 580645 703156
rect 579843 702948 579909 702949
rect 579843 702884 579844 702948
rect 579908 702884 579909 702948
rect 579843 702883 579909 702884
rect 579659 702404 579725 702405
rect 579659 702340 579660 702404
rect 579724 702340 579725 702404
rect 579659 702339 579725 702340
rect 579662 696557 579722 702339
rect 579846 697645 579906 702883
rect 580027 700908 580093 700909
rect 580027 700844 580028 700908
rect 580092 700844 580093 700908
rect 580027 700843 580093 700844
rect 579843 697644 579909 697645
rect 579843 697580 579844 697644
rect 579908 697580 579909 697644
rect 579843 697579 579909 697580
rect 579659 696556 579725 696557
rect 579659 696492 579660 696556
rect 579724 696492 579725 696556
rect 579659 696491 579725 696492
rect 580030 683909 580090 700843
rect 580395 700772 580461 700773
rect 580395 700708 580396 700772
rect 580460 700708 580461 700772
rect 580395 700707 580461 700708
rect 580211 700636 580277 700637
rect 580211 700572 580212 700636
rect 580276 700572 580277 700636
rect 580211 700571 580277 700572
rect 580214 697237 580274 700571
rect 580211 697236 580277 697237
rect 580211 697172 580212 697236
rect 580276 697172 580277 697236
rect 580211 697171 580277 697172
rect 580398 696690 580458 700707
rect 580214 696630 580458 696690
rect 580027 683908 580093 683909
rect 580027 683844 580028 683908
rect 580092 683844 580093 683908
rect 580027 683843 580093 683844
rect 577638 634770 578066 634830
rect 578006 617541 578066 634770
rect 578003 617540 578069 617541
rect 578003 617476 578004 617540
rect 578068 617476 578069 617540
rect 578003 617475 578069 617476
rect 577454 576810 578066 576870
rect 578006 564365 578066 576810
rect 578003 564364 578069 564365
rect 578003 564300 578004 564364
rect 578068 564300 578069 564364
rect 578003 564299 578069 564300
rect 580214 458149 580274 696630
rect 580395 696556 580461 696557
rect 580395 696492 580396 696556
rect 580460 696492 580461 696556
rect 580395 696491 580461 696492
rect 580398 511325 580458 696491
rect 580582 591021 580642 703155
rect 582419 701996 582485 701997
rect 582419 701932 582420 701996
rect 582484 701932 582485 701996
rect 582419 701931 582485 701932
rect 580947 701180 581013 701181
rect 580947 701116 580948 701180
rect 581012 701116 581013 701180
rect 580947 701115 581013 701116
rect 580763 697644 580829 697645
rect 580763 697580 580764 697644
rect 580828 697580 580829 697644
rect 580763 697579 580829 697580
rect 580766 670717 580826 697579
rect 580763 670716 580829 670717
rect 580763 670652 580764 670716
rect 580828 670652 580829 670716
rect 580763 670651 580829 670652
rect 580579 591020 580645 591021
rect 580579 590956 580580 591020
rect 580644 590956 580645 591020
rect 580579 590955 580645 590956
rect 580950 579597 581010 701115
rect 580947 579596 581013 579597
rect 580947 579532 580948 579596
rect 581012 579532 581013 579596
rect 580947 579531 581013 579532
rect 580395 511324 580461 511325
rect 580395 511260 580396 511324
rect 580460 511260 580461 511324
rect 580395 511259 580461 511260
rect 580211 458148 580277 458149
rect 580211 458084 580212 458148
rect 580276 458084 580277 458148
rect 580211 458083 580277 458084
rect 577270 364290 578066 364350
rect 578006 351933 578066 364290
rect 578003 351932 578069 351933
rect 578003 351868 578004 351932
rect 578068 351868 578069 351932
rect 578003 351867 578069 351868
rect 577794 291454 578414 301784
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 572667 33148 572733 33149
rect 572667 33084 572668 33148
rect 572732 33084 572733 33148
rect 572667 33083 572733 33084
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 295174 582134 299784
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 582422 179213 582482 701931
rect 582603 699956 582669 699957
rect 582603 699892 582604 699956
rect 582668 699892 582669 699956
rect 582603 699891 582669 699892
rect 582606 192541 582666 699891
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 582603 192540 582669 192541
rect 582603 192476 582604 192540
rect 582668 192476 582669 192540
rect 582603 192475 582669 192476
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 582419 179212 582485 179213
rect 582419 179148 582420 179212
rect 582484 179148 582485 179212
rect 582419 179147 582485 179148
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 187034 687218 187270 687454
rect 187034 686898 187270 687134
rect 202394 669218 202630 669454
rect 202394 668898 202630 669134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 187034 651218 187270 651454
rect 187034 650898 187270 651134
rect 202394 633218 202630 633454
rect 202394 632898 202630 633134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 187034 615218 187270 615454
rect 187034 614898 187270 615134
rect 202394 597218 202630 597454
rect 202394 596898 202630 597134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 187034 579218 187270 579454
rect 187034 578898 187270 579134
rect 202394 561218 202630 561454
rect 202394 560898 202630 561134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 187034 543218 187270 543454
rect 187034 542898 187270 543134
rect 202394 525218 202630 525454
rect 202394 524898 202630 525134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 187034 507218 187270 507454
rect 187034 506898 187270 507134
rect 202394 489218 202630 489454
rect 202394 488898 202630 489134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 187034 471218 187270 471454
rect 187034 470898 187270 471134
rect 202394 453218 202630 453454
rect 202394 452898 202630 453134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 187034 435218 187270 435454
rect 187034 434898 187270 435134
rect 202394 417218 202630 417454
rect 202394 416898 202630 417134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 187034 399218 187270 399454
rect 187034 398898 187270 399134
rect 202394 381218 202630 381454
rect 202394 380898 202630 381134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 187034 363218 187270 363454
rect 187034 362898 187270 363134
rect 202394 345218 202630 345454
rect 202394 344898 202630 345134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 187034 327218 187270 327454
rect 187034 326898 187270 327134
rect 202394 309218 202630 309454
rect 202394 308898 202630 309134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 217754 687218 217990 687454
rect 217754 686898 217990 687134
rect 217754 651218 217990 651454
rect 217754 650898 217990 651134
rect 217754 615218 217990 615454
rect 217754 614898 217990 615134
rect 217754 579218 217990 579454
rect 217754 578898 217990 579134
rect 217754 543218 217990 543454
rect 217754 542898 217990 543134
rect 217754 507218 217990 507454
rect 217754 506898 217990 507134
rect 217754 471218 217990 471454
rect 217754 470898 217990 471134
rect 217754 435218 217990 435454
rect 217754 434898 217990 435134
rect 217754 399218 217990 399454
rect 217754 398898 217990 399134
rect 217754 363218 217990 363454
rect 217754 362898 217990 363134
rect 217754 327218 217990 327454
rect 217754 326898 217990 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 248474 687218 248710 687454
rect 248474 686898 248710 687134
rect 279194 687218 279430 687454
rect 279194 686898 279430 687134
rect 309914 687218 310150 687454
rect 309914 686898 310150 687134
rect 340634 687218 340870 687454
rect 340634 686898 340870 687134
rect 371354 687218 371590 687454
rect 371354 686898 371590 687134
rect 402074 687218 402310 687454
rect 402074 686898 402310 687134
rect 432794 687218 433030 687454
rect 432794 686898 433030 687134
rect 463514 687218 463750 687454
rect 463514 686898 463750 687134
rect 494234 687218 494470 687454
rect 494234 686898 494470 687134
rect 233114 669218 233350 669454
rect 233114 668898 233350 669134
rect 263834 669218 264070 669454
rect 263834 668898 264070 669134
rect 294554 669218 294790 669454
rect 294554 668898 294790 669134
rect 325274 669218 325510 669454
rect 325274 668898 325510 669134
rect 355994 669218 356230 669454
rect 355994 668898 356230 669134
rect 386714 669218 386950 669454
rect 386714 668898 386950 669134
rect 417434 669218 417670 669454
rect 417434 668898 417670 669134
rect 448154 669218 448390 669454
rect 448154 668898 448390 669134
rect 478874 669218 479110 669454
rect 478874 668898 479110 669134
rect 509594 669218 509830 669454
rect 509594 668898 509830 669134
rect 248474 651218 248710 651454
rect 248474 650898 248710 651134
rect 279194 651218 279430 651454
rect 279194 650898 279430 651134
rect 309914 651218 310150 651454
rect 309914 650898 310150 651134
rect 340634 651218 340870 651454
rect 340634 650898 340870 651134
rect 371354 651218 371590 651454
rect 371354 650898 371590 651134
rect 402074 651218 402310 651454
rect 402074 650898 402310 651134
rect 432794 651218 433030 651454
rect 432794 650898 433030 651134
rect 463514 651218 463750 651454
rect 463514 650898 463750 651134
rect 494234 651218 494470 651454
rect 494234 650898 494470 651134
rect 233114 633218 233350 633454
rect 233114 632898 233350 633134
rect 263834 633218 264070 633454
rect 263834 632898 264070 633134
rect 294554 633218 294790 633454
rect 294554 632898 294790 633134
rect 325274 633218 325510 633454
rect 325274 632898 325510 633134
rect 355994 633218 356230 633454
rect 355994 632898 356230 633134
rect 386714 633218 386950 633454
rect 386714 632898 386950 633134
rect 417434 633218 417670 633454
rect 417434 632898 417670 633134
rect 448154 633218 448390 633454
rect 448154 632898 448390 633134
rect 478874 633218 479110 633454
rect 478874 632898 479110 633134
rect 509594 633218 509830 633454
rect 509594 632898 509830 633134
rect 248474 615218 248710 615454
rect 248474 614898 248710 615134
rect 279194 615218 279430 615454
rect 279194 614898 279430 615134
rect 309914 615218 310150 615454
rect 309914 614898 310150 615134
rect 340634 615218 340870 615454
rect 340634 614898 340870 615134
rect 371354 615218 371590 615454
rect 371354 614898 371590 615134
rect 402074 615218 402310 615454
rect 402074 614898 402310 615134
rect 432794 615218 433030 615454
rect 432794 614898 433030 615134
rect 463514 615218 463750 615454
rect 463514 614898 463750 615134
rect 494234 615218 494470 615454
rect 494234 614898 494470 615134
rect 233114 597218 233350 597454
rect 233114 596898 233350 597134
rect 263834 597218 264070 597454
rect 263834 596898 264070 597134
rect 294554 597218 294790 597454
rect 294554 596898 294790 597134
rect 325274 597218 325510 597454
rect 325274 596898 325510 597134
rect 355994 597218 356230 597454
rect 355994 596898 356230 597134
rect 386714 597218 386950 597454
rect 386714 596898 386950 597134
rect 417434 597218 417670 597454
rect 417434 596898 417670 597134
rect 448154 597218 448390 597454
rect 448154 596898 448390 597134
rect 478874 597218 479110 597454
rect 478874 596898 479110 597134
rect 509594 597218 509830 597454
rect 509594 596898 509830 597134
rect 248474 579218 248710 579454
rect 248474 578898 248710 579134
rect 279194 579218 279430 579454
rect 279194 578898 279430 579134
rect 309914 579218 310150 579454
rect 309914 578898 310150 579134
rect 340634 579218 340870 579454
rect 340634 578898 340870 579134
rect 371354 579218 371590 579454
rect 371354 578898 371590 579134
rect 402074 579218 402310 579454
rect 402074 578898 402310 579134
rect 432794 579218 433030 579454
rect 432794 578898 433030 579134
rect 463514 579218 463750 579454
rect 463514 578898 463750 579134
rect 494234 579218 494470 579454
rect 494234 578898 494470 579134
rect 233114 561218 233350 561454
rect 233114 560898 233350 561134
rect 263834 561218 264070 561454
rect 263834 560898 264070 561134
rect 294554 561218 294790 561454
rect 294554 560898 294790 561134
rect 325274 561218 325510 561454
rect 325274 560898 325510 561134
rect 355994 561218 356230 561454
rect 355994 560898 356230 561134
rect 386714 561218 386950 561454
rect 386714 560898 386950 561134
rect 417434 561218 417670 561454
rect 417434 560898 417670 561134
rect 448154 561218 448390 561454
rect 448154 560898 448390 561134
rect 478874 561218 479110 561454
rect 478874 560898 479110 561134
rect 509594 561218 509830 561454
rect 509594 560898 509830 561134
rect 248474 543218 248710 543454
rect 248474 542898 248710 543134
rect 279194 543218 279430 543454
rect 279194 542898 279430 543134
rect 309914 543218 310150 543454
rect 309914 542898 310150 543134
rect 340634 543218 340870 543454
rect 340634 542898 340870 543134
rect 371354 543218 371590 543454
rect 371354 542898 371590 543134
rect 402074 543218 402310 543454
rect 402074 542898 402310 543134
rect 432794 543218 433030 543454
rect 432794 542898 433030 543134
rect 463514 543218 463750 543454
rect 463514 542898 463750 543134
rect 494234 543218 494470 543454
rect 494234 542898 494470 543134
rect 233114 525218 233350 525454
rect 233114 524898 233350 525134
rect 263834 525218 264070 525454
rect 263834 524898 264070 525134
rect 294554 525218 294790 525454
rect 294554 524898 294790 525134
rect 325274 525218 325510 525454
rect 325274 524898 325510 525134
rect 355994 525218 356230 525454
rect 355994 524898 356230 525134
rect 386714 525218 386950 525454
rect 386714 524898 386950 525134
rect 417434 525218 417670 525454
rect 417434 524898 417670 525134
rect 448154 525218 448390 525454
rect 448154 524898 448390 525134
rect 478874 525218 479110 525454
rect 478874 524898 479110 525134
rect 509594 525218 509830 525454
rect 509594 524898 509830 525134
rect 248474 507218 248710 507454
rect 248474 506898 248710 507134
rect 279194 507218 279430 507454
rect 279194 506898 279430 507134
rect 309914 507218 310150 507454
rect 309914 506898 310150 507134
rect 340634 507218 340870 507454
rect 340634 506898 340870 507134
rect 371354 507218 371590 507454
rect 371354 506898 371590 507134
rect 402074 507218 402310 507454
rect 402074 506898 402310 507134
rect 432794 507218 433030 507454
rect 432794 506898 433030 507134
rect 463514 507218 463750 507454
rect 463514 506898 463750 507134
rect 494234 507218 494470 507454
rect 494234 506898 494470 507134
rect 233114 489218 233350 489454
rect 233114 488898 233350 489134
rect 263834 489218 264070 489454
rect 263834 488898 264070 489134
rect 294554 489218 294790 489454
rect 294554 488898 294790 489134
rect 325274 489218 325510 489454
rect 325274 488898 325510 489134
rect 355994 489218 356230 489454
rect 355994 488898 356230 489134
rect 386714 489218 386950 489454
rect 386714 488898 386950 489134
rect 417434 489218 417670 489454
rect 417434 488898 417670 489134
rect 448154 489218 448390 489454
rect 448154 488898 448390 489134
rect 478874 489218 479110 489454
rect 478874 488898 479110 489134
rect 509594 489218 509830 489454
rect 509594 488898 509830 489134
rect 248474 471218 248710 471454
rect 248474 470898 248710 471134
rect 279194 471218 279430 471454
rect 279194 470898 279430 471134
rect 309914 471218 310150 471454
rect 309914 470898 310150 471134
rect 340634 471218 340870 471454
rect 340634 470898 340870 471134
rect 371354 471218 371590 471454
rect 371354 470898 371590 471134
rect 402074 471218 402310 471454
rect 402074 470898 402310 471134
rect 432794 471218 433030 471454
rect 432794 470898 433030 471134
rect 463514 471218 463750 471454
rect 463514 470898 463750 471134
rect 494234 471218 494470 471454
rect 494234 470898 494470 471134
rect 233114 453218 233350 453454
rect 233114 452898 233350 453134
rect 263834 453218 264070 453454
rect 263834 452898 264070 453134
rect 294554 453218 294790 453454
rect 294554 452898 294790 453134
rect 325274 453218 325510 453454
rect 325274 452898 325510 453134
rect 355994 453218 356230 453454
rect 355994 452898 356230 453134
rect 386714 453218 386950 453454
rect 386714 452898 386950 453134
rect 417434 453218 417670 453454
rect 417434 452898 417670 453134
rect 448154 453218 448390 453454
rect 448154 452898 448390 453134
rect 478874 453218 479110 453454
rect 478874 452898 479110 453134
rect 509594 453218 509830 453454
rect 509594 452898 509830 453134
rect 248474 435218 248710 435454
rect 248474 434898 248710 435134
rect 279194 435218 279430 435454
rect 279194 434898 279430 435134
rect 309914 435218 310150 435454
rect 309914 434898 310150 435134
rect 340634 435218 340870 435454
rect 340634 434898 340870 435134
rect 371354 435218 371590 435454
rect 371354 434898 371590 435134
rect 402074 435218 402310 435454
rect 402074 434898 402310 435134
rect 432794 435218 433030 435454
rect 432794 434898 433030 435134
rect 463514 435218 463750 435454
rect 463514 434898 463750 435134
rect 494234 435218 494470 435454
rect 494234 434898 494470 435134
rect 233114 417218 233350 417454
rect 233114 416898 233350 417134
rect 263834 417218 264070 417454
rect 263834 416898 264070 417134
rect 294554 417218 294790 417454
rect 294554 416898 294790 417134
rect 325274 417218 325510 417454
rect 325274 416898 325510 417134
rect 355994 417218 356230 417454
rect 355994 416898 356230 417134
rect 386714 417218 386950 417454
rect 386714 416898 386950 417134
rect 417434 417218 417670 417454
rect 417434 416898 417670 417134
rect 448154 417218 448390 417454
rect 448154 416898 448390 417134
rect 478874 417218 479110 417454
rect 478874 416898 479110 417134
rect 509594 417218 509830 417454
rect 509594 416898 509830 417134
rect 248474 399218 248710 399454
rect 248474 398898 248710 399134
rect 279194 399218 279430 399454
rect 279194 398898 279430 399134
rect 309914 399218 310150 399454
rect 309914 398898 310150 399134
rect 340634 399218 340870 399454
rect 340634 398898 340870 399134
rect 371354 399218 371590 399454
rect 371354 398898 371590 399134
rect 402074 399218 402310 399454
rect 402074 398898 402310 399134
rect 432794 399218 433030 399454
rect 432794 398898 433030 399134
rect 463514 399218 463750 399454
rect 463514 398898 463750 399134
rect 494234 399218 494470 399454
rect 494234 398898 494470 399134
rect 233114 381218 233350 381454
rect 233114 380898 233350 381134
rect 263834 381218 264070 381454
rect 263834 380898 264070 381134
rect 294554 381218 294790 381454
rect 294554 380898 294790 381134
rect 325274 381218 325510 381454
rect 325274 380898 325510 381134
rect 355994 381218 356230 381454
rect 355994 380898 356230 381134
rect 386714 381218 386950 381454
rect 386714 380898 386950 381134
rect 417434 381218 417670 381454
rect 417434 380898 417670 381134
rect 448154 381218 448390 381454
rect 448154 380898 448390 381134
rect 478874 381218 479110 381454
rect 478874 380898 479110 381134
rect 509594 381218 509830 381454
rect 509594 380898 509830 381134
rect 248474 363218 248710 363454
rect 248474 362898 248710 363134
rect 279194 363218 279430 363454
rect 279194 362898 279430 363134
rect 309914 363218 310150 363454
rect 309914 362898 310150 363134
rect 340634 363218 340870 363454
rect 340634 362898 340870 363134
rect 371354 363218 371590 363454
rect 371354 362898 371590 363134
rect 402074 363218 402310 363454
rect 402074 362898 402310 363134
rect 432794 363218 433030 363454
rect 432794 362898 433030 363134
rect 463514 363218 463750 363454
rect 463514 362898 463750 363134
rect 494234 363218 494470 363454
rect 494234 362898 494470 363134
rect 233114 345218 233350 345454
rect 233114 344898 233350 345134
rect 263834 345218 264070 345454
rect 263834 344898 264070 345134
rect 294554 345218 294790 345454
rect 294554 344898 294790 345134
rect 325274 345218 325510 345454
rect 325274 344898 325510 345134
rect 355994 345218 356230 345454
rect 355994 344898 356230 345134
rect 386714 345218 386950 345454
rect 386714 344898 386950 345134
rect 417434 345218 417670 345454
rect 417434 344898 417670 345134
rect 448154 345218 448390 345454
rect 448154 344898 448390 345134
rect 478874 345218 479110 345454
rect 478874 344898 479110 345134
rect 509594 345218 509830 345454
rect 509594 344898 509830 345134
rect 248474 327218 248710 327454
rect 248474 326898 248710 327134
rect 279194 327218 279430 327454
rect 279194 326898 279430 327134
rect 309914 327218 310150 327454
rect 309914 326898 310150 327134
rect 340634 327218 340870 327454
rect 340634 326898 340870 327134
rect 371354 327218 371590 327454
rect 371354 326898 371590 327134
rect 402074 327218 402310 327454
rect 402074 326898 402310 327134
rect 432794 327218 433030 327454
rect 432794 326898 433030 327134
rect 463514 327218 463750 327454
rect 463514 326898 463750 327134
rect 494234 327218 494470 327454
rect 494234 326898 494470 327134
rect 233114 309218 233350 309454
rect 233114 308898 233350 309134
rect 263834 309218 264070 309454
rect 263834 308898 264070 309134
rect 294554 309218 294790 309454
rect 294554 308898 294790 309134
rect 325274 309218 325510 309454
rect 325274 308898 325510 309134
rect 355994 309218 356230 309454
rect 355994 308898 356230 309134
rect 386714 309218 386950 309454
rect 386714 308898 386950 309134
rect 417434 309218 417670 309454
rect 417434 308898 417670 309134
rect 448154 309218 448390 309454
rect 448154 308898 448390 309134
rect 478874 309218 479110 309454
rect 478874 308898 479110 309134
rect 509594 309218 509830 309454
rect 509594 308898 509830 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 524954 687218 525190 687454
rect 524954 686898 525190 687134
rect 524954 651218 525190 651454
rect 524954 650898 525190 651134
rect 524954 615218 525190 615454
rect 524954 614898 525190 615134
rect 524954 579218 525190 579454
rect 524954 578898 525190 579134
rect 524954 543218 525190 543454
rect 524954 542898 525190 543134
rect 524954 507218 525190 507454
rect 524954 506898 525190 507134
rect 524954 471218 525190 471454
rect 524954 470898 525190 471134
rect 524954 435218 525190 435454
rect 524954 434898 525190 435134
rect 524954 399218 525190 399454
rect 524954 398898 525190 399134
rect 524954 363218 525190 363454
rect 524954 362898 525190 363134
rect 524954 327218 525190 327454
rect 524954 326898 525190 327134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 540314 669218 540550 669454
rect 540314 668898 540550 669134
rect 540314 633218 540550 633454
rect 540314 632898 540550 633134
rect 540314 597218 540550 597454
rect 540314 596898 540550 597134
rect 540314 561218 540550 561454
rect 540314 560898 540550 561134
rect 540314 525218 540550 525454
rect 540314 524898 540550 525134
rect 540314 489218 540550 489454
rect 540314 488898 540550 489134
rect 540314 453218 540550 453454
rect 540314 452898 540550 453134
rect 540314 417218 540550 417454
rect 540314 416898 540550 417134
rect 540314 381218 540550 381454
rect 540314 380898 540550 381134
rect 540314 345218 540550 345454
rect 540314 344898 540550 345134
rect 540314 309218 540550 309454
rect 540314 308898 540550 309134
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 555674 687218 555910 687454
rect 555674 686898 555910 687134
rect 555674 651218 555910 651454
rect 555674 650898 555910 651134
rect 555674 615218 555910 615454
rect 555674 614898 555910 615134
rect 555674 579218 555910 579454
rect 555674 578898 555910 579134
rect 555674 543218 555910 543454
rect 555674 542898 555910 543134
rect 555674 507218 555910 507454
rect 555674 506898 555910 507134
rect 555674 471218 555910 471454
rect 555674 470898 555910 471134
rect 555674 435218 555910 435454
rect 555674 434898 555910 435134
rect 555674 399218 555910 399454
rect 555674 398898 555910 399134
rect 555674 363218 555910 363454
rect 555674 362898 555910 363134
rect 555674 327218 555910 327454
rect 555674 326898 555910 327134
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 571034 669218 571270 669454
rect 571034 668898 571270 669134
rect 571034 633218 571270 633454
rect 571034 632898 571270 633134
rect 571034 597218 571270 597454
rect 571034 596898 571270 597134
rect 571034 561218 571270 561454
rect 571034 560898 571270 561134
rect 571034 525218 571270 525454
rect 571034 524898 571270 525134
rect 571034 489218 571270 489454
rect 571034 488898 571270 489134
rect 571034 453218 571270 453454
rect 571034 452898 571270 453134
rect 571034 417218 571270 417454
rect 571034 416898 571270 417134
rect 571034 381218 571270 381454
rect 571034 380898 571270 381134
rect 571034 345218 571270 345454
rect 571034 344898 571270 345134
rect 571034 309218 571270 309454
rect 571034 308898 571270 309134
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 187034 687454
rect 187270 687218 217754 687454
rect 217990 687218 248474 687454
rect 248710 687218 279194 687454
rect 279430 687218 309914 687454
rect 310150 687218 340634 687454
rect 340870 687218 371354 687454
rect 371590 687218 402074 687454
rect 402310 687218 432794 687454
rect 433030 687218 463514 687454
rect 463750 687218 494234 687454
rect 494470 687218 524954 687454
rect 525190 687218 555674 687454
rect 555910 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 187034 687134
rect 187270 686898 217754 687134
rect 217990 686898 248474 687134
rect 248710 686898 279194 687134
rect 279430 686898 309914 687134
rect 310150 686898 340634 687134
rect 340870 686898 371354 687134
rect 371590 686898 402074 687134
rect 402310 686898 432794 687134
rect 433030 686898 463514 687134
rect 463750 686898 494234 687134
rect 494470 686898 524954 687134
rect 525190 686898 555674 687134
rect 555910 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 202394 669454
rect 202630 669218 233114 669454
rect 233350 669218 263834 669454
rect 264070 669218 294554 669454
rect 294790 669218 325274 669454
rect 325510 669218 355994 669454
rect 356230 669218 386714 669454
rect 386950 669218 417434 669454
rect 417670 669218 448154 669454
rect 448390 669218 478874 669454
rect 479110 669218 509594 669454
rect 509830 669218 540314 669454
rect 540550 669218 571034 669454
rect 571270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 202394 669134
rect 202630 668898 233114 669134
rect 233350 668898 263834 669134
rect 264070 668898 294554 669134
rect 294790 668898 325274 669134
rect 325510 668898 355994 669134
rect 356230 668898 386714 669134
rect 386950 668898 417434 669134
rect 417670 668898 448154 669134
rect 448390 668898 478874 669134
rect 479110 668898 509594 669134
rect 509830 668898 540314 669134
rect 540550 668898 571034 669134
rect 571270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 187034 651454
rect 187270 651218 217754 651454
rect 217990 651218 248474 651454
rect 248710 651218 279194 651454
rect 279430 651218 309914 651454
rect 310150 651218 340634 651454
rect 340870 651218 371354 651454
rect 371590 651218 402074 651454
rect 402310 651218 432794 651454
rect 433030 651218 463514 651454
rect 463750 651218 494234 651454
rect 494470 651218 524954 651454
rect 525190 651218 555674 651454
rect 555910 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 187034 651134
rect 187270 650898 217754 651134
rect 217990 650898 248474 651134
rect 248710 650898 279194 651134
rect 279430 650898 309914 651134
rect 310150 650898 340634 651134
rect 340870 650898 371354 651134
rect 371590 650898 402074 651134
rect 402310 650898 432794 651134
rect 433030 650898 463514 651134
rect 463750 650898 494234 651134
rect 494470 650898 524954 651134
rect 525190 650898 555674 651134
rect 555910 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 202394 633454
rect 202630 633218 233114 633454
rect 233350 633218 263834 633454
rect 264070 633218 294554 633454
rect 294790 633218 325274 633454
rect 325510 633218 355994 633454
rect 356230 633218 386714 633454
rect 386950 633218 417434 633454
rect 417670 633218 448154 633454
rect 448390 633218 478874 633454
rect 479110 633218 509594 633454
rect 509830 633218 540314 633454
rect 540550 633218 571034 633454
rect 571270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 202394 633134
rect 202630 632898 233114 633134
rect 233350 632898 263834 633134
rect 264070 632898 294554 633134
rect 294790 632898 325274 633134
rect 325510 632898 355994 633134
rect 356230 632898 386714 633134
rect 386950 632898 417434 633134
rect 417670 632898 448154 633134
rect 448390 632898 478874 633134
rect 479110 632898 509594 633134
rect 509830 632898 540314 633134
rect 540550 632898 571034 633134
rect 571270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 187034 615454
rect 187270 615218 217754 615454
rect 217990 615218 248474 615454
rect 248710 615218 279194 615454
rect 279430 615218 309914 615454
rect 310150 615218 340634 615454
rect 340870 615218 371354 615454
rect 371590 615218 402074 615454
rect 402310 615218 432794 615454
rect 433030 615218 463514 615454
rect 463750 615218 494234 615454
rect 494470 615218 524954 615454
rect 525190 615218 555674 615454
rect 555910 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 187034 615134
rect 187270 614898 217754 615134
rect 217990 614898 248474 615134
rect 248710 614898 279194 615134
rect 279430 614898 309914 615134
rect 310150 614898 340634 615134
rect 340870 614898 371354 615134
rect 371590 614898 402074 615134
rect 402310 614898 432794 615134
rect 433030 614898 463514 615134
rect 463750 614898 494234 615134
rect 494470 614898 524954 615134
rect 525190 614898 555674 615134
rect 555910 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 202394 597454
rect 202630 597218 233114 597454
rect 233350 597218 263834 597454
rect 264070 597218 294554 597454
rect 294790 597218 325274 597454
rect 325510 597218 355994 597454
rect 356230 597218 386714 597454
rect 386950 597218 417434 597454
rect 417670 597218 448154 597454
rect 448390 597218 478874 597454
rect 479110 597218 509594 597454
rect 509830 597218 540314 597454
rect 540550 597218 571034 597454
rect 571270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 202394 597134
rect 202630 596898 233114 597134
rect 233350 596898 263834 597134
rect 264070 596898 294554 597134
rect 294790 596898 325274 597134
rect 325510 596898 355994 597134
rect 356230 596898 386714 597134
rect 386950 596898 417434 597134
rect 417670 596898 448154 597134
rect 448390 596898 478874 597134
rect 479110 596898 509594 597134
rect 509830 596898 540314 597134
rect 540550 596898 571034 597134
rect 571270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 187034 579454
rect 187270 579218 217754 579454
rect 217990 579218 248474 579454
rect 248710 579218 279194 579454
rect 279430 579218 309914 579454
rect 310150 579218 340634 579454
rect 340870 579218 371354 579454
rect 371590 579218 402074 579454
rect 402310 579218 432794 579454
rect 433030 579218 463514 579454
rect 463750 579218 494234 579454
rect 494470 579218 524954 579454
rect 525190 579218 555674 579454
rect 555910 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 187034 579134
rect 187270 578898 217754 579134
rect 217990 578898 248474 579134
rect 248710 578898 279194 579134
rect 279430 578898 309914 579134
rect 310150 578898 340634 579134
rect 340870 578898 371354 579134
rect 371590 578898 402074 579134
rect 402310 578898 432794 579134
rect 433030 578898 463514 579134
rect 463750 578898 494234 579134
rect 494470 578898 524954 579134
rect 525190 578898 555674 579134
rect 555910 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 202394 561454
rect 202630 561218 233114 561454
rect 233350 561218 263834 561454
rect 264070 561218 294554 561454
rect 294790 561218 325274 561454
rect 325510 561218 355994 561454
rect 356230 561218 386714 561454
rect 386950 561218 417434 561454
rect 417670 561218 448154 561454
rect 448390 561218 478874 561454
rect 479110 561218 509594 561454
rect 509830 561218 540314 561454
rect 540550 561218 571034 561454
rect 571270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 202394 561134
rect 202630 560898 233114 561134
rect 233350 560898 263834 561134
rect 264070 560898 294554 561134
rect 294790 560898 325274 561134
rect 325510 560898 355994 561134
rect 356230 560898 386714 561134
rect 386950 560898 417434 561134
rect 417670 560898 448154 561134
rect 448390 560898 478874 561134
rect 479110 560898 509594 561134
rect 509830 560898 540314 561134
rect 540550 560898 571034 561134
rect 571270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 187034 543454
rect 187270 543218 217754 543454
rect 217990 543218 248474 543454
rect 248710 543218 279194 543454
rect 279430 543218 309914 543454
rect 310150 543218 340634 543454
rect 340870 543218 371354 543454
rect 371590 543218 402074 543454
rect 402310 543218 432794 543454
rect 433030 543218 463514 543454
rect 463750 543218 494234 543454
rect 494470 543218 524954 543454
rect 525190 543218 555674 543454
rect 555910 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 187034 543134
rect 187270 542898 217754 543134
rect 217990 542898 248474 543134
rect 248710 542898 279194 543134
rect 279430 542898 309914 543134
rect 310150 542898 340634 543134
rect 340870 542898 371354 543134
rect 371590 542898 402074 543134
rect 402310 542898 432794 543134
rect 433030 542898 463514 543134
rect 463750 542898 494234 543134
rect 494470 542898 524954 543134
rect 525190 542898 555674 543134
rect 555910 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 202394 525454
rect 202630 525218 233114 525454
rect 233350 525218 263834 525454
rect 264070 525218 294554 525454
rect 294790 525218 325274 525454
rect 325510 525218 355994 525454
rect 356230 525218 386714 525454
rect 386950 525218 417434 525454
rect 417670 525218 448154 525454
rect 448390 525218 478874 525454
rect 479110 525218 509594 525454
rect 509830 525218 540314 525454
rect 540550 525218 571034 525454
rect 571270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 202394 525134
rect 202630 524898 233114 525134
rect 233350 524898 263834 525134
rect 264070 524898 294554 525134
rect 294790 524898 325274 525134
rect 325510 524898 355994 525134
rect 356230 524898 386714 525134
rect 386950 524898 417434 525134
rect 417670 524898 448154 525134
rect 448390 524898 478874 525134
rect 479110 524898 509594 525134
rect 509830 524898 540314 525134
rect 540550 524898 571034 525134
rect 571270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 187034 507454
rect 187270 507218 217754 507454
rect 217990 507218 248474 507454
rect 248710 507218 279194 507454
rect 279430 507218 309914 507454
rect 310150 507218 340634 507454
rect 340870 507218 371354 507454
rect 371590 507218 402074 507454
rect 402310 507218 432794 507454
rect 433030 507218 463514 507454
rect 463750 507218 494234 507454
rect 494470 507218 524954 507454
rect 525190 507218 555674 507454
rect 555910 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 187034 507134
rect 187270 506898 217754 507134
rect 217990 506898 248474 507134
rect 248710 506898 279194 507134
rect 279430 506898 309914 507134
rect 310150 506898 340634 507134
rect 340870 506898 371354 507134
rect 371590 506898 402074 507134
rect 402310 506898 432794 507134
rect 433030 506898 463514 507134
rect 463750 506898 494234 507134
rect 494470 506898 524954 507134
rect 525190 506898 555674 507134
rect 555910 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 202394 489454
rect 202630 489218 233114 489454
rect 233350 489218 263834 489454
rect 264070 489218 294554 489454
rect 294790 489218 325274 489454
rect 325510 489218 355994 489454
rect 356230 489218 386714 489454
rect 386950 489218 417434 489454
rect 417670 489218 448154 489454
rect 448390 489218 478874 489454
rect 479110 489218 509594 489454
rect 509830 489218 540314 489454
rect 540550 489218 571034 489454
rect 571270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 202394 489134
rect 202630 488898 233114 489134
rect 233350 488898 263834 489134
rect 264070 488898 294554 489134
rect 294790 488898 325274 489134
rect 325510 488898 355994 489134
rect 356230 488898 386714 489134
rect 386950 488898 417434 489134
rect 417670 488898 448154 489134
rect 448390 488898 478874 489134
rect 479110 488898 509594 489134
rect 509830 488898 540314 489134
rect 540550 488898 571034 489134
rect 571270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 187034 471454
rect 187270 471218 217754 471454
rect 217990 471218 248474 471454
rect 248710 471218 279194 471454
rect 279430 471218 309914 471454
rect 310150 471218 340634 471454
rect 340870 471218 371354 471454
rect 371590 471218 402074 471454
rect 402310 471218 432794 471454
rect 433030 471218 463514 471454
rect 463750 471218 494234 471454
rect 494470 471218 524954 471454
rect 525190 471218 555674 471454
rect 555910 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 187034 471134
rect 187270 470898 217754 471134
rect 217990 470898 248474 471134
rect 248710 470898 279194 471134
rect 279430 470898 309914 471134
rect 310150 470898 340634 471134
rect 340870 470898 371354 471134
rect 371590 470898 402074 471134
rect 402310 470898 432794 471134
rect 433030 470898 463514 471134
rect 463750 470898 494234 471134
rect 494470 470898 524954 471134
rect 525190 470898 555674 471134
rect 555910 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 202394 453454
rect 202630 453218 233114 453454
rect 233350 453218 263834 453454
rect 264070 453218 294554 453454
rect 294790 453218 325274 453454
rect 325510 453218 355994 453454
rect 356230 453218 386714 453454
rect 386950 453218 417434 453454
rect 417670 453218 448154 453454
rect 448390 453218 478874 453454
rect 479110 453218 509594 453454
rect 509830 453218 540314 453454
rect 540550 453218 571034 453454
rect 571270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 202394 453134
rect 202630 452898 233114 453134
rect 233350 452898 263834 453134
rect 264070 452898 294554 453134
rect 294790 452898 325274 453134
rect 325510 452898 355994 453134
rect 356230 452898 386714 453134
rect 386950 452898 417434 453134
rect 417670 452898 448154 453134
rect 448390 452898 478874 453134
rect 479110 452898 509594 453134
rect 509830 452898 540314 453134
rect 540550 452898 571034 453134
rect 571270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 187034 435454
rect 187270 435218 217754 435454
rect 217990 435218 248474 435454
rect 248710 435218 279194 435454
rect 279430 435218 309914 435454
rect 310150 435218 340634 435454
rect 340870 435218 371354 435454
rect 371590 435218 402074 435454
rect 402310 435218 432794 435454
rect 433030 435218 463514 435454
rect 463750 435218 494234 435454
rect 494470 435218 524954 435454
rect 525190 435218 555674 435454
rect 555910 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 187034 435134
rect 187270 434898 217754 435134
rect 217990 434898 248474 435134
rect 248710 434898 279194 435134
rect 279430 434898 309914 435134
rect 310150 434898 340634 435134
rect 340870 434898 371354 435134
rect 371590 434898 402074 435134
rect 402310 434898 432794 435134
rect 433030 434898 463514 435134
rect 463750 434898 494234 435134
rect 494470 434898 524954 435134
rect 525190 434898 555674 435134
rect 555910 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 202394 417454
rect 202630 417218 233114 417454
rect 233350 417218 263834 417454
rect 264070 417218 294554 417454
rect 294790 417218 325274 417454
rect 325510 417218 355994 417454
rect 356230 417218 386714 417454
rect 386950 417218 417434 417454
rect 417670 417218 448154 417454
rect 448390 417218 478874 417454
rect 479110 417218 509594 417454
rect 509830 417218 540314 417454
rect 540550 417218 571034 417454
rect 571270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 202394 417134
rect 202630 416898 233114 417134
rect 233350 416898 263834 417134
rect 264070 416898 294554 417134
rect 294790 416898 325274 417134
rect 325510 416898 355994 417134
rect 356230 416898 386714 417134
rect 386950 416898 417434 417134
rect 417670 416898 448154 417134
rect 448390 416898 478874 417134
rect 479110 416898 509594 417134
rect 509830 416898 540314 417134
rect 540550 416898 571034 417134
rect 571270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 187034 399454
rect 187270 399218 217754 399454
rect 217990 399218 248474 399454
rect 248710 399218 279194 399454
rect 279430 399218 309914 399454
rect 310150 399218 340634 399454
rect 340870 399218 371354 399454
rect 371590 399218 402074 399454
rect 402310 399218 432794 399454
rect 433030 399218 463514 399454
rect 463750 399218 494234 399454
rect 494470 399218 524954 399454
rect 525190 399218 555674 399454
rect 555910 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 187034 399134
rect 187270 398898 217754 399134
rect 217990 398898 248474 399134
rect 248710 398898 279194 399134
rect 279430 398898 309914 399134
rect 310150 398898 340634 399134
rect 340870 398898 371354 399134
rect 371590 398898 402074 399134
rect 402310 398898 432794 399134
rect 433030 398898 463514 399134
rect 463750 398898 494234 399134
rect 494470 398898 524954 399134
rect 525190 398898 555674 399134
rect 555910 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 202394 381454
rect 202630 381218 233114 381454
rect 233350 381218 263834 381454
rect 264070 381218 294554 381454
rect 294790 381218 325274 381454
rect 325510 381218 355994 381454
rect 356230 381218 386714 381454
rect 386950 381218 417434 381454
rect 417670 381218 448154 381454
rect 448390 381218 478874 381454
rect 479110 381218 509594 381454
rect 509830 381218 540314 381454
rect 540550 381218 571034 381454
rect 571270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 202394 381134
rect 202630 380898 233114 381134
rect 233350 380898 263834 381134
rect 264070 380898 294554 381134
rect 294790 380898 325274 381134
rect 325510 380898 355994 381134
rect 356230 380898 386714 381134
rect 386950 380898 417434 381134
rect 417670 380898 448154 381134
rect 448390 380898 478874 381134
rect 479110 380898 509594 381134
rect 509830 380898 540314 381134
rect 540550 380898 571034 381134
rect 571270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 187034 363454
rect 187270 363218 217754 363454
rect 217990 363218 248474 363454
rect 248710 363218 279194 363454
rect 279430 363218 309914 363454
rect 310150 363218 340634 363454
rect 340870 363218 371354 363454
rect 371590 363218 402074 363454
rect 402310 363218 432794 363454
rect 433030 363218 463514 363454
rect 463750 363218 494234 363454
rect 494470 363218 524954 363454
rect 525190 363218 555674 363454
rect 555910 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 187034 363134
rect 187270 362898 217754 363134
rect 217990 362898 248474 363134
rect 248710 362898 279194 363134
rect 279430 362898 309914 363134
rect 310150 362898 340634 363134
rect 340870 362898 371354 363134
rect 371590 362898 402074 363134
rect 402310 362898 432794 363134
rect 433030 362898 463514 363134
rect 463750 362898 494234 363134
rect 494470 362898 524954 363134
rect 525190 362898 555674 363134
rect 555910 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 202394 345454
rect 202630 345218 233114 345454
rect 233350 345218 263834 345454
rect 264070 345218 294554 345454
rect 294790 345218 325274 345454
rect 325510 345218 355994 345454
rect 356230 345218 386714 345454
rect 386950 345218 417434 345454
rect 417670 345218 448154 345454
rect 448390 345218 478874 345454
rect 479110 345218 509594 345454
rect 509830 345218 540314 345454
rect 540550 345218 571034 345454
rect 571270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 202394 345134
rect 202630 344898 233114 345134
rect 233350 344898 263834 345134
rect 264070 344898 294554 345134
rect 294790 344898 325274 345134
rect 325510 344898 355994 345134
rect 356230 344898 386714 345134
rect 386950 344898 417434 345134
rect 417670 344898 448154 345134
rect 448390 344898 478874 345134
rect 479110 344898 509594 345134
rect 509830 344898 540314 345134
rect 540550 344898 571034 345134
rect 571270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 187034 327454
rect 187270 327218 217754 327454
rect 217990 327218 248474 327454
rect 248710 327218 279194 327454
rect 279430 327218 309914 327454
rect 310150 327218 340634 327454
rect 340870 327218 371354 327454
rect 371590 327218 402074 327454
rect 402310 327218 432794 327454
rect 433030 327218 463514 327454
rect 463750 327218 494234 327454
rect 494470 327218 524954 327454
rect 525190 327218 555674 327454
rect 555910 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 187034 327134
rect 187270 326898 217754 327134
rect 217990 326898 248474 327134
rect 248710 326898 279194 327134
rect 279430 326898 309914 327134
rect 310150 326898 340634 327134
rect 340870 326898 371354 327134
rect 371590 326898 402074 327134
rect 402310 326898 432794 327134
rect 433030 326898 463514 327134
rect 463750 326898 494234 327134
rect 494470 326898 524954 327134
rect 525190 326898 555674 327134
rect 555910 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 202394 309454
rect 202630 309218 233114 309454
rect 233350 309218 263834 309454
rect 264070 309218 294554 309454
rect 294790 309218 325274 309454
rect 325510 309218 355994 309454
rect 356230 309218 386714 309454
rect 386950 309218 417434 309454
rect 417670 309218 448154 309454
rect 448390 309218 478874 309454
rect 479110 309218 509594 309454
rect 509830 309218 540314 309454
rect 540550 309218 571034 309454
rect 571270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 202394 309134
rect 202630 308898 233114 309134
rect 233350 308898 263834 309134
rect 264070 308898 294554 309134
rect 294790 308898 325274 309134
rect 325510 308898 355994 309134
rect 356230 308898 386714 309134
rect 386950 308898 417434 309134
rect 417670 308898 448154 309134
rect 448390 308898 478874 309134
rect 479110 308898 509594 309134
rect 509830 308898 540314 309134
rect 540550 308898 571034 309134
rect 571270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use computer  computer
timestamp 1634795968
transform 1 0 182784 0 1 301784
box 381 0 399634 400000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 301784 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 701784 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 701784 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 701784 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 701784 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 701784 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 701784 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 701784 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 701784 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 701784 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 701784 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 701784 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 299784 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 703784 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 703784 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 703784 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 703784 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 703784 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 703784 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 703784 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 703784 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 703784 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 703784 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 703784 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 703784 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 299784 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 703784 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 703784 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 703784 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 703784 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 703784 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 703784 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 703784 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 703784 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 703784 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 703784 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 703784 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 299784 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 703784 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 703784 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 703784 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 703784 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 703784 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 703784 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 703784 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 703784 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 703784 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 703784 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 703784 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 299784 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 703784 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 703784 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 703784 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 703784 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 703784 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 703784 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 703784 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 703784 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 703784 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 703784 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 703784 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 299784 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 703784 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 703784 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 703784 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 703784 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 703784 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 703784 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 703784 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 703784 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 703784 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 703784 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 703784 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 301784 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 701784 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 701784 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 701784 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 701784 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 701784 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 701784 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 701784 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 701784 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 701784 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 701784 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 701784 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 299784 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 703784 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 703784 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 703784 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 703784 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 703784 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 703784 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 703784 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 703784 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 703784 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 703784 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 703784 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
