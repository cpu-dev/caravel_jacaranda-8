VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO computer
  CLASS BLOCK ;
  FOREIGN computer ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 996.000 4.510 1000.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 996.000 267.630 1000.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 996.000 293.850 1000.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 996.000 320.070 1000.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 996.000 346.290 1000.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 996.000 372.510 1000.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 996.000 399.190 1000.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 996.000 425.410 1000.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 996.000 451.630 1000.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 996.000 477.850 1000.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 996.000 504.530 1000.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 996.000 30.730 1000.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 996.000 530.750 1000.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 996.000 556.970 1000.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 996.000 583.190 1000.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 996.000 609.410 1000.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 996.000 636.090 1000.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 996.000 662.310 1000.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 996.000 688.530 1000.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 996.000 714.750 1000.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 996.000 740.970 1000.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 996.000 767.650 1000.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 996.000 56.950 1000.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 996.000 793.870 1000.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 996.000 820.090 1000.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 996.000 846.310 1000.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 996.000 872.530 1000.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 996.000 899.210 1000.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.150 996.000 925.430 1000.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 996.000 951.650 1000.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.590 996.000 977.870 1000.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 996.000 83.170 1000.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 996.000 109.390 1000.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 996.000 136.070 1000.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 996.000 162.290 1000.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 996.000 188.510 1000.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 996.000 214.730 1000.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 996.000 240.950 1000.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 996.000 13.250 1000.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 996.000 276.370 1000.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 996.000 302.590 1000.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 996.000 328.810 1000.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 996.000 355.030 1000.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 996.000 381.710 1000.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 996.000 407.930 1000.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 996.000 434.150 1000.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 996.000 460.370 1000.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 996.000 486.590 1000.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 996.000 513.270 1000.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 996.000 39.470 1000.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 996.000 539.490 1000.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 996.000 565.710 1000.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 996.000 591.930 1000.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 996.000 618.150 1000.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 996.000 644.830 1000.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 996.000 671.050 1000.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 996.000 697.270 1000.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 996.000 723.490 1000.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 996.000 749.710 1000.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 996.000 776.390 1000.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 996.000 65.690 1000.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 996.000 802.610 1000.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 996.000 828.830 1000.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 996.000 855.050 1000.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 996.000 881.730 1000.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.670 996.000 907.950 1000.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 996.000 934.170 1000.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 996.000 960.390 1000.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330 996.000 986.610 1000.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 996.000 91.910 1000.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 996.000 118.130 1000.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 996.000 144.810 1000.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 996.000 171.030 1000.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 996.000 197.250 1000.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 996.000 223.470 1000.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 996.000 249.690 1000.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 996.000 21.990 1000.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 996.000 285.110 1000.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 996.000 311.330 1000.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 996.000 337.550 1000.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 996.000 363.770 1000.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 996.000 390.450 1000.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 996.000 416.670 1000.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 996.000 442.890 1000.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 996.000 469.110 1000.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 996.000 495.330 1000.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 996.000 522.010 1000.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 996.000 48.210 1000.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 996.000 548.230 1000.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 996.000 574.450 1000.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 996.000 600.670 1000.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 996.000 626.890 1000.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 996.000 653.570 1000.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 996.000 679.790 1000.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 996.000 706.010 1000.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 996.000 732.230 1000.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.630 996.000 758.910 1000.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 996.000 785.130 1000.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 996.000 74.430 1000.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 996.000 811.350 1000.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 996.000 837.570 1000.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 996.000 863.790 1000.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 996.000 890.470 1000.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 996.000 916.690 1000.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 996.000 942.910 1000.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 996.000 969.130 1000.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 996.000 995.350 1000.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 996.000 100.650 1000.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 996.000 126.870 1000.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 996.000 153.550 1000.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 996.000 179.770 1000.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 996.000 205.990 1000.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 996.000 232.210 1000.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 996.000 258.890 1000.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.610 0.000 994.890 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 0.000 997.190 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 0.000 830.670 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 0.000 836.650 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.810 0.000 843.090 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 0.000 867.010 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 0.000 873.450 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 0.000 885.410 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 0.000 891.390 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 0.000 903.810 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.490 0.000 915.770 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 0.000 922.210 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 0.000 928.190 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.870 0.000 940.150 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.850 0.000 946.130 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 0.000 952.570 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.270 0.000 958.550 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.250 0.000 964.530 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 0.000 970.510 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 0.000 976.950 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 0.000 611.710 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 0.000 642.070 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 0.000 648.050 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 0.000 672.430 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 0.000 684.850 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 0.000 696.810 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 0.000 739.590 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 0.000 751.550 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 0.000 781.910 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 0.000 787.890 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 0.000 812.270 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.230 0.000 832.510 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 0.000 844.930 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 0.000 850.910 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 0.000 869.310 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 0.000 887.710 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 0.000 893.690 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 0.000 905.650 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 0.000 924.050 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 0.000 930.030 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 0.000 936.010 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 0.000 948.430 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 0.000 954.410 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 0.000 960.390 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 0.000 966.830 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.510 0.000 978.790 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.490 0.000 984.770 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 0.000 990.750 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 0.000 510.050 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 0.000 662.310 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 0.000 735.450 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 0.000 759.830 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 0.000 765.810 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 0.000 784.210 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 0.000 820.550 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 0.000 846.770 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 0.000 859.190 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 0.000 865.170 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 0.000 877.590 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 0.000 883.570 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 0.000 889.550 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.670 0.000 907.950 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.630 0.000 919.910 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 0.000 925.890 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 0.000 938.310 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 0.000 956.250 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 0.000 962.690 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 0.000 968.670 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.370 0.000 974.650 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 0.000 987.070 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.770 0.000 993.050 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 0.000 597.450 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 0.000 609.410 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 0.000 694.970 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 0.000 712.910 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 0.000 743.270 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 0.000 774.090 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 0.000 792.030 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 0.000 798.470 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 0.000 816.410 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 987.600 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.060 987.445 ;
      LAYER met1 ;
        RECT 2.830 8.540 999.050 987.600 ;
      LAYER met2 ;
        RECT 0.090 995.720 3.950 996.000 ;
        RECT 4.790 995.720 12.690 996.000 ;
        RECT 13.530 995.720 21.430 996.000 ;
        RECT 22.270 995.720 30.170 996.000 ;
        RECT 31.010 995.720 38.910 996.000 ;
        RECT 39.750 995.720 47.650 996.000 ;
        RECT 48.490 995.720 56.390 996.000 ;
        RECT 57.230 995.720 65.130 996.000 ;
        RECT 65.970 995.720 73.870 996.000 ;
        RECT 74.710 995.720 82.610 996.000 ;
        RECT 83.450 995.720 91.350 996.000 ;
        RECT 92.190 995.720 100.090 996.000 ;
        RECT 100.930 995.720 108.830 996.000 ;
        RECT 109.670 995.720 117.570 996.000 ;
        RECT 118.410 995.720 126.310 996.000 ;
        RECT 127.150 995.720 135.510 996.000 ;
        RECT 136.350 995.720 144.250 996.000 ;
        RECT 145.090 995.720 152.990 996.000 ;
        RECT 153.830 995.720 161.730 996.000 ;
        RECT 162.570 995.720 170.470 996.000 ;
        RECT 171.310 995.720 179.210 996.000 ;
        RECT 180.050 995.720 187.950 996.000 ;
        RECT 188.790 995.720 196.690 996.000 ;
        RECT 197.530 995.720 205.430 996.000 ;
        RECT 206.270 995.720 214.170 996.000 ;
        RECT 215.010 995.720 222.910 996.000 ;
        RECT 223.750 995.720 231.650 996.000 ;
        RECT 232.490 995.720 240.390 996.000 ;
        RECT 241.230 995.720 249.130 996.000 ;
        RECT 249.970 995.720 258.330 996.000 ;
        RECT 259.170 995.720 267.070 996.000 ;
        RECT 267.910 995.720 275.810 996.000 ;
        RECT 276.650 995.720 284.550 996.000 ;
        RECT 285.390 995.720 293.290 996.000 ;
        RECT 294.130 995.720 302.030 996.000 ;
        RECT 302.870 995.720 310.770 996.000 ;
        RECT 311.610 995.720 319.510 996.000 ;
        RECT 320.350 995.720 328.250 996.000 ;
        RECT 329.090 995.720 336.990 996.000 ;
        RECT 337.830 995.720 345.730 996.000 ;
        RECT 346.570 995.720 354.470 996.000 ;
        RECT 355.310 995.720 363.210 996.000 ;
        RECT 364.050 995.720 371.950 996.000 ;
        RECT 372.790 995.720 381.150 996.000 ;
        RECT 381.990 995.720 389.890 996.000 ;
        RECT 390.730 995.720 398.630 996.000 ;
        RECT 399.470 995.720 407.370 996.000 ;
        RECT 408.210 995.720 416.110 996.000 ;
        RECT 416.950 995.720 424.850 996.000 ;
        RECT 425.690 995.720 433.590 996.000 ;
        RECT 434.430 995.720 442.330 996.000 ;
        RECT 443.170 995.720 451.070 996.000 ;
        RECT 451.910 995.720 459.810 996.000 ;
        RECT 460.650 995.720 468.550 996.000 ;
        RECT 469.390 995.720 477.290 996.000 ;
        RECT 478.130 995.720 486.030 996.000 ;
        RECT 486.870 995.720 494.770 996.000 ;
        RECT 495.610 995.720 503.970 996.000 ;
        RECT 504.810 995.720 512.710 996.000 ;
        RECT 513.550 995.720 521.450 996.000 ;
        RECT 522.290 995.720 530.190 996.000 ;
        RECT 531.030 995.720 538.930 996.000 ;
        RECT 539.770 995.720 547.670 996.000 ;
        RECT 548.510 995.720 556.410 996.000 ;
        RECT 557.250 995.720 565.150 996.000 ;
        RECT 565.990 995.720 573.890 996.000 ;
        RECT 574.730 995.720 582.630 996.000 ;
        RECT 583.470 995.720 591.370 996.000 ;
        RECT 592.210 995.720 600.110 996.000 ;
        RECT 600.950 995.720 608.850 996.000 ;
        RECT 609.690 995.720 617.590 996.000 ;
        RECT 618.430 995.720 626.330 996.000 ;
        RECT 627.170 995.720 635.530 996.000 ;
        RECT 636.370 995.720 644.270 996.000 ;
        RECT 645.110 995.720 653.010 996.000 ;
        RECT 653.850 995.720 661.750 996.000 ;
        RECT 662.590 995.720 670.490 996.000 ;
        RECT 671.330 995.720 679.230 996.000 ;
        RECT 680.070 995.720 687.970 996.000 ;
        RECT 688.810 995.720 696.710 996.000 ;
        RECT 697.550 995.720 705.450 996.000 ;
        RECT 706.290 995.720 714.190 996.000 ;
        RECT 715.030 995.720 722.930 996.000 ;
        RECT 723.770 995.720 731.670 996.000 ;
        RECT 732.510 995.720 740.410 996.000 ;
        RECT 741.250 995.720 749.150 996.000 ;
        RECT 749.990 995.720 758.350 996.000 ;
        RECT 759.190 995.720 767.090 996.000 ;
        RECT 767.930 995.720 775.830 996.000 ;
        RECT 776.670 995.720 784.570 996.000 ;
        RECT 785.410 995.720 793.310 996.000 ;
        RECT 794.150 995.720 802.050 996.000 ;
        RECT 802.890 995.720 810.790 996.000 ;
        RECT 811.630 995.720 819.530 996.000 ;
        RECT 820.370 995.720 828.270 996.000 ;
        RECT 829.110 995.720 837.010 996.000 ;
        RECT 837.850 995.720 845.750 996.000 ;
        RECT 846.590 995.720 854.490 996.000 ;
        RECT 855.330 995.720 863.230 996.000 ;
        RECT 864.070 995.720 871.970 996.000 ;
        RECT 872.810 995.720 881.170 996.000 ;
        RECT 882.010 995.720 889.910 996.000 ;
        RECT 890.750 995.720 898.650 996.000 ;
        RECT 899.490 995.720 907.390 996.000 ;
        RECT 908.230 995.720 916.130 996.000 ;
        RECT 916.970 995.720 924.870 996.000 ;
        RECT 925.710 995.720 933.610 996.000 ;
        RECT 934.450 995.720 942.350 996.000 ;
        RECT 943.190 995.720 951.090 996.000 ;
        RECT 951.930 995.720 959.830 996.000 ;
        RECT 960.670 995.720 968.570 996.000 ;
        RECT 969.410 995.720 977.310 996.000 ;
        RECT 978.150 995.720 986.050 996.000 ;
        RECT 986.890 995.720 994.790 996.000 ;
        RECT 995.630 995.720 999.020 996.000 ;
        RECT 0.090 4.280 999.020 995.720 ;
        RECT 0.090 3.670 0.730 4.280 ;
        RECT 1.570 3.670 2.570 4.280 ;
        RECT 3.410 3.670 4.410 4.280 ;
        RECT 5.250 3.670 6.710 4.280 ;
        RECT 7.550 3.670 8.550 4.280 ;
        RECT 9.390 3.670 10.850 4.280 ;
        RECT 11.690 3.670 12.690 4.280 ;
        RECT 13.530 3.670 14.530 4.280 ;
        RECT 15.370 3.670 16.830 4.280 ;
        RECT 17.670 3.670 18.670 4.280 ;
        RECT 19.510 3.670 20.970 4.280 ;
        RECT 21.810 3.670 22.810 4.280 ;
        RECT 23.650 3.670 24.650 4.280 ;
        RECT 25.490 3.670 26.950 4.280 ;
        RECT 27.790 3.670 28.790 4.280 ;
        RECT 29.630 3.670 31.090 4.280 ;
        RECT 31.930 3.670 32.930 4.280 ;
        RECT 33.770 3.670 34.770 4.280 ;
        RECT 35.610 3.670 37.070 4.280 ;
        RECT 37.910 3.670 38.910 4.280 ;
        RECT 39.750 3.670 41.210 4.280 ;
        RECT 42.050 3.670 43.050 4.280 ;
        RECT 43.890 3.670 45.350 4.280 ;
        RECT 46.190 3.670 47.190 4.280 ;
        RECT 48.030 3.670 49.030 4.280 ;
        RECT 49.870 3.670 51.330 4.280 ;
        RECT 52.170 3.670 53.170 4.280 ;
        RECT 54.010 3.670 55.470 4.280 ;
        RECT 56.310 3.670 57.310 4.280 ;
        RECT 58.150 3.670 59.150 4.280 ;
        RECT 59.990 3.670 61.450 4.280 ;
        RECT 62.290 3.670 63.290 4.280 ;
        RECT 64.130 3.670 65.590 4.280 ;
        RECT 66.430 3.670 67.430 4.280 ;
        RECT 68.270 3.670 69.270 4.280 ;
        RECT 70.110 3.670 71.570 4.280 ;
        RECT 72.410 3.670 73.410 4.280 ;
        RECT 74.250 3.670 75.710 4.280 ;
        RECT 76.550 3.670 77.550 4.280 ;
        RECT 78.390 3.670 79.390 4.280 ;
        RECT 80.230 3.670 81.690 4.280 ;
        RECT 82.530 3.670 83.530 4.280 ;
        RECT 84.370 3.670 85.830 4.280 ;
        RECT 86.670 3.670 87.670 4.280 ;
        RECT 88.510 3.670 89.970 4.280 ;
        RECT 90.810 3.670 91.810 4.280 ;
        RECT 92.650 3.670 93.650 4.280 ;
        RECT 94.490 3.670 95.950 4.280 ;
        RECT 96.790 3.670 97.790 4.280 ;
        RECT 98.630 3.670 100.090 4.280 ;
        RECT 100.930 3.670 101.930 4.280 ;
        RECT 102.770 3.670 103.770 4.280 ;
        RECT 104.610 3.670 106.070 4.280 ;
        RECT 106.910 3.670 107.910 4.280 ;
        RECT 108.750 3.670 110.210 4.280 ;
        RECT 111.050 3.670 112.050 4.280 ;
        RECT 112.890 3.670 113.890 4.280 ;
        RECT 114.730 3.670 116.190 4.280 ;
        RECT 117.030 3.670 118.030 4.280 ;
        RECT 118.870 3.670 120.330 4.280 ;
        RECT 121.170 3.670 122.170 4.280 ;
        RECT 123.010 3.670 124.010 4.280 ;
        RECT 124.850 3.670 126.310 4.280 ;
        RECT 127.150 3.670 128.150 4.280 ;
        RECT 128.990 3.670 130.450 4.280 ;
        RECT 131.290 3.670 132.290 4.280 ;
        RECT 133.130 3.670 134.590 4.280 ;
        RECT 135.430 3.670 136.430 4.280 ;
        RECT 137.270 3.670 138.270 4.280 ;
        RECT 139.110 3.670 140.570 4.280 ;
        RECT 141.410 3.670 142.410 4.280 ;
        RECT 143.250 3.670 144.710 4.280 ;
        RECT 145.550 3.670 146.550 4.280 ;
        RECT 147.390 3.670 148.390 4.280 ;
        RECT 149.230 3.670 150.690 4.280 ;
        RECT 151.530 3.670 152.530 4.280 ;
        RECT 153.370 3.670 154.830 4.280 ;
        RECT 155.670 3.670 156.670 4.280 ;
        RECT 157.510 3.670 158.510 4.280 ;
        RECT 159.350 3.670 160.810 4.280 ;
        RECT 161.650 3.670 162.650 4.280 ;
        RECT 163.490 3.670 164.950 4.280 ;
        RECT 165.790 3.670 166.790 4.280 ;
        RECT 167.630 3.670 169.090 4.280 ;
        RECT 169.930 3.670 170.930 4.280 ;
        RECT 171.770 3.670 172.770 4.280 ;
        RECT 173.610 3.670 175.070 4.280 ;
        RECT 175.910 3.670 176.910 4.280 ;
        RECT 177.750 3.670 179.210 4.280 ;
        RECT 180.050 3.670 181.050 4.280 ;
        RECT 181.890 3.670 182.890 4.280 ;
        RECT 183.730 3.670 185.190 4.280 ;
        RECT 186.030 3.670 187.030 4.280 ;
        RECT 187.870 3.670 189.330 4.280 ;
        RECT 190.170 3.670 191.170 4.280 ;
        RECT 192.010 3.670 193.010 4.280 ;
        RECT 193.850 3.670 195.310 4.280 ;
        RECT 196.150 3.670 197.150 4.280 ;
        RECT 197.990 3.670 199.450 4.280 ;
        RECT 200.290 3.670 201.290 4.280 ;
        RECT 202.130 3.670 203.130 4.280 ;
        RECT 203.970 3.670 205.430 4.280 ;
        RECT 206.270 3.670 207.270 4.280 ;
        RECT 208.110 3.670 209.570 4.280 ;
        RECT 210.410 3.670 211.410 4.280 ;
        RECT 212.250 3.670 213.710 4.280 ;
        RECT 214.550 3.670 215.550 4.280 ;
        RECT 216.390 3.670 217.390 4.280 ;
        RECT 218.230 3.670 219.690 4.280 ;
        RECT 220.530 3.670 221.530 4.280 ;
        RECT 222.370 3.670 223.830 4.280 ;
        RECT 224.670 3.670 225.670 4.280 ;
        RECT 226.510 3.670 227.510 4.280 ;
        RECT 228.350 3.670 229.810 4.280 ;
        RECT 230.650 3.670 231.650 4.280 ;
        RECT 232.490 3.670 233.950 4.280 ;
        RECT 234.790 3.670 235.790 4.280 ;
        RECT 236.630 3.670 237.630 4.280 ;
        RECT 238.470 3.670 239.930 4.280 ;
        RECT 240.770 3.670 241.770 4.280 ;
        RECT 242.610 3.670 244.070 4.280 ;
        RECT 244.910 3.670 245.910 4.280 ;
        RECT 246.750 3.670 247.750 4.280 ;
        RECT 248.590 3.670 250.050 4.280 ;
        RECT 250.890 3.670 251.890 4.280 ;
        RECT 252.730 3.670 254.190 4.280 ;
        RECT 255.030 3.670 256.030 4.280 ;
        RECT 256.870 3.670 258.330 4.280 ;
        RECT 259.170 3.670 260.170 4.280 ;
        RECT 261.010 3.670 262.010 4.280 ;
        RECT 262.850 3.670 264.310 4.280 ;
        RECT 265.150 3.670 266.150 4.280 ;
        RECT 266.990 3.670 268.450 4.280 ;
        RECT 269.290 3.670 270.290 4.280 ;
        RECT 271.130 3.670 272.130 4.280 ;
        RECT 272.970 3.670 274.430 4.280 ;
        RECT 275.270 3.670 276.270 4.280 ;
        RECT 277.110 3.670 278.570 4.280 ;
        RECT 279.410 3.670 280.410 4.280 ;
        RECT 281.250 3.670 282.250 4.280 ;
        RECT 283.090 3.670 284.550 4.280 ;
        RECT 285.390 3.670 286.390 4.280 ;
        RECT 287.230 3.670 288.690 4.280 ;
        RECT 289.530 3.670 290.530 4.280 ;
        RECT 291.370 3.670 292.830 4.280 ;
        RECT 293.670 3.670 294.670 4.280 ;
        RECT 295.510 3.670 296.510 4.280 ;
        RECT 297.350 3.670 298.810 4.280 ;
        RECT 299.650 3.670 300.650 4.280 ;
        RECT 301.490 3.670 302.950 4.280 ;
        RECT 303.790 3.670 304.790 4.280 ;
        RECT 305.630 3.670 306.630 4.280 ;
        RECT 307.470 3.670 308.930 4.280 ;
        RECT 309.770 3.670 310.770 4.280 ;
        RECT 311.610 3.670 313.070 4.280 ;
        RECT 313.910 3.670 314.910 4.280 ;
        RECT 315.750 3.670 316.750 4.280 ;
        RECT 317.590 3.670 319.050 4.280 ;
        RECT 319.890 3.670 320.890 4.280 ;
        RECT 321.730 3.670 323.190 4.280 ;
        RECT 324.030 3.670 325.030 4.280 ;
        RECT 325.870 3.670 326.870 4.280 ;
        RECT 327.710 3.670 329.170 4.280 ;
        RECT 330.010 3.670 331.010 4.280 ;
        RECT 331.850 3.670 333.310 4.280 ;
        RECT 334.150 3.670 335.150 4.280 ;
        RECT 335.990 3.670 337.450 4.280 ;
        RECT 338.290 3.670 339.290 4.280 ;
        RECT 340.130 3.670 341.130 4.280 ;
        RECT 341.970 3.670 343.430 4.280 ;
        RECT 344.270 3.670 345.270 4.280 ;
        RECT 346.110 3.670 347.570 4.280 ;
        RECT 348.410 3.670 349.410 4.280 ;
        RECT 350.250 3.670 351.250 4.280 ;
        RECT 352.090 3.670 353.550 4.280 ;
        RECT 354.390 3.670 355.390 4.280 ;
        RECT 356.230 3.670 357.690 4.280 ;
        RECT 358.530 3.670 359.530 4.280 ;
        RECT 360.370 3.670 361.370 4.280 ;
        RECT 362.210 3.670 363.670 4.280 ;
        RECT 364.510 3.670 365.510 4.280 ;
        RECT 366.350 3.670 367.810 4.280 ;
        RECT 368.650 3.670 369.650 4.280 ;
        RECT 370.490 3.670 371.490 4.280 ;
        RECT 372.330 3.670 373.790 4.280 ;
        RECT 374.630 3.670 375.630 4.280 ;
        RECT 376.470 3.670 377.930 4.280 ;
        RECT 378.770 3.670 379.770 4.280 ;
        RECT 380.610 3.670 382.070 4.280 ;
        RECT 382.910 3.670 383.910 4.280 ;
        RECT 384.750 3.670 385.750 4.280 ;
        RECT 386.590 3.670 388.050 4.280 ;
        RECT 388.890 3.670 389.890 4.280 ;
        RECT 390.730 3.670 392.190 4.280 ;
        RECT 393.030 3.670 394.030 4.280 ;
        RECT 394.870 3.670 395.870 4.280 ;
        RECT 396.710 3.670 398.170 4.280 ;
        RECT 399.010 3.670 400.010 4.280 ;
        RECT 400.850 3.670 402.310 4.280 ;
        RECT 403.150 3.670 404.150 4.280 ;
        RECT 404.990 3.670 405.990 4.280 ;
        RECT 406.830 3.670 408.290 4.280 ;
        RECT 409.130 3.670 410.130 4.280 ;
        RECT 410.970 3.670 412.430 4.280 ;
        RECT 413.270 3.670 414.270 4.280 ;
        RECT 415.110 3.670 416.110 4.280 ;
        RECT 416.950 3.670 418.410 4.280 ;
        RECT 419.250 3.670 420.250 4.280 ;
        RECT 421.090 3.670 422.550 4.280 ;
        RECT 423.390 3.670 424.390 4.280 ;
        RECT 425.230 3.670 426.690 4.280 ;
        RECT 427.530 3.670 428.530 4.280 ;
        RECT 429.370 3.670 430.370 4.280 ;
        RECT 431.210 3.670 432.670 4.280 ;
        RECT 433.510 3.670 434.510 4.280 ;
        RECT 435.350 3.670 436.810 4.280 ;
        RECT 437.650 3.670 438.650 4.280 ;
        RECT 439.490 3.670 440.490 4.280 ;
        RECT 441.330 3.670 442.790 4.280 ;
        RECT 443.630 3.670 444.630 4.280 ;
        RECT 445.470 3.670 446.930 4.280 ;
        RECT 447.770 3.670 448.770 4.280 ;
        RECT 449.610 3.670 450.610 4.280 ;
        RECT 451.450 3.670 452.910 4.280 ;
        RECT 453.750 3.670 454.750 4.280 ;
        RECT 455.590 3.670 457.050 4.280 ;
        RECT 457.890 3.670 458.890 4.280 ;
        RECT 459.730 3.670 461.190 4.280 ;
        RECT 462.030 3.670 463.030 4.280 ;
        RECT 463.870 3.670 464.870 4.280 ;
        RECT 465.710 3.670 467.170 4.280 ;
        RECT 468.010 3.670 469.010 4.280 ;
        RECT 469.850 3.670 471.310 4.280 ;
        RECT 472.150 3.670 473.150 4.280 ;
        RECT 473.990 3.670 474.990 4.280 ;
        RECT 475.830 3.670 477.290 4.280 ;
        RECT 478.130 3.670 479.130 4.280 ;
        RECT 479.970 3.670 481.430 4.280 ;
        RECT 482.270 3.670 483.270 4.280 ;
        RECT 484.110 3.670 485.110 4.280 ;
        RECT 485.950 3.670 487.410 4.280 ;
        RECT 488.250 3.670 489.250 4.280 ;
        RECT 490.090 3.670 491.550 4.280 ;
        RECT 492.390 3.670 493.390 4.280 ;
        RECT 494.230 3.670 495.230 4.280 ;
        RECT 496.070 3.670 497.530 4.280 ;
        RECT 498.370 3.670 499.370 4.280 ;
        RECT 500.210 3.670 501.670 4.280 ;
        RECT 502.510 3.670 503.510 4.280 ;
        RECT 504.350 3.670 505.810 4.280 ;
        RECT 506.650 3.670 507.650 4.280 ;
        RECT 508.490 3.670 509.490 4.280 ;
        RECT 510.330 3.670 511.790 4.280 ;
        RECT 512.630 3.670 513.630 4.280 ;
        RECT 514.470 3.670 515.930 4.280 ;
        RECT 516.770 3.670 517.770 4.280 ;
        RECT 518.610 3.670 519.610 4.280 ;
        RECT 520.450 3.670 521.910 4.280 ;
        RECT 522.750 3.670 523.750 4.280 ;
        RECT 524.590 3.670 526.050 4.280 ;
        RECT 526.890 3.670 527.890 4.280 ;
        RECT 528.730 3.670 529.730 4.280 ;
        RECT 530.570 3.670 532.030 4.280 ;
        RECT 532.870 3.670 533.870 4.280 ;
        RECT 534.710 3.670 536.170 4.280 ;
        RECT 537.010 3.670 538.010 4.280 ;
        RECT 538.850 3.670 539.850 4.280 ;
        RECT 540.690 3.670 542.150 4.280 ;
        RECT 542.990 3.670 543.990 4.280 ;
        RECT 544.830 3.670 546.290 4.280 ;
        RECT 547.130 3.670 548.130 4.280 ;
        RECT 548.970 3.670 550.430 4.280 ;
        RECT 551.270 3.670 552.270 4.280 ;
        RECT 553.110 3.670 554.110 4.280 ;
        RECT 554.950 3.670 556.410 4.280 ;
        RECT 557.250 3.670 558.250 4.280 ;
        RECT 559.090 3.670 560.550 4.280 ;
        RECT 561.390 3.670 562.390 4.280 ;
        RECT 563.230 3.670 564.230 4.280 ;
        RECT 565.070 3.670 566.530 4.280 ;
        RECT 567.370 3.670 568.370 4.280 ;
        RECT 569.210 3.670 570.670 4.280 ;
        RECT 571.510 3.670 572.510 4.280 ;
        RECT 573.350 3.670 574.350 4.280 ;
        RECT 575.190 3.670 576.650 4.280 ;
        RECT 577.490 3.670 578.490 4.280 ;
        RECT 579.330 3.670 580.790 4.280 ;
        RECT 581.630 3.670 582.630 4.280 ;
        RECT 583.470 3.670 584.930 4.280 ;
        RECT 585.770 3.670 586.770 4.280 ;
        RECT 587.610 3.670 588.610 4.280 ;
        RECT 589.450 3.670 590.910 4.280 ;
        RECT 591.750 3.670 592.750 4.280 ;
        RECT 593.590 3.670 595.050 4.280 ;
        RECT 595.890 3.670 596.890 4.280 ;
        RECT 597.730 3.670 598.730 4.280 ;
        RECT 599.570 3.670 601.030 4.280 ;
        RECT 601.870 3.670 602.870 4.280 ;
        RECT 603.710 3.670 605.170 4.280 ;
        RECT 606.010 3.670 607.010 4.280 ;
        RECT 607.850 3.670 608.850 4.280 ;
        RECT 609.690 3.670 611.150 4.280 ;
        RECT 611.990 3.670 612.990 4.280 ;
        RECT 613.830 3.670 615.290 4.280 ;
        RECT 616.130 3.670 617.130 4.280 ;
        RECT 617.970 3.670 618.970 4.280 ;
        RECT 619.810 3.670 621.270 4.280 ;
        RECT 622.110 3.670 623.110 4.280 ;
        RECT 623.950 3.670 625.410 4.280 ;
        RECT 626.250 3.670 627.250 4.280 ;
        RECT 628.090 3.670 629.550 4.280 ;
        RECT 630.390 3.670 631.390 4.280 ;
        RECT 632.230 3.670 633.230 4.280 ;
        RECT 634.070 3.670 635.530 4.280 ;
        RECT 636.370 3.670 637.370 4.280 ;
        RECT 638.210 3.670 639.670 4.280 ;
        RECT 640.510 3.670 641.510 4.280 ;
        RECT 642.350 3.670 643.350 4.280 ;
        RECT 644.190 3.670 645.650 4.280 ;
        RECT 646.490 3.670 647.490 4.280 ;
        RECT 648.330 3.670 649.790 4.280 ;
        RECT 650.630 3.670 651.630 4.280 ;
        RECT 652.470 3.670 653.470 4.280 ;
        RECT 654.310 3.670 655.770 4.280 ;
        RECT 656.610 3.670 657.610 4.280 ;
        RECT 658.450 3.670 659.910 4.280 ;
        RECT 660.750 3.670 661.750 4.280 ;
        RECT 662.590 3.670 663.590 4.280 ;
        RECT 664.430 3.670 665.890 4.280 ;
        RECT 666.730 3.670 667.730 4.280 ;
        RECT 668.570 3.670 670.030 4.280 ;
        RECT 670.870 3.670 671.870 4.280 ;
        RECT 672.710 3.670 674.170 4.280 ;
        RECT 675.010 3.670 676.010 4.280 ;
        RECT 676.850 3.670 677.850 4.280 ;
        RECT 678.690 3.670 680.150 4.280 ;
        RECT 680.990 3.670 681.990 4.280 ;
        RECT 682.830 3.670 684.290 4.280 ;
        RECT 685.130 3.670 686.130 4.280 ;
        RECT 686.970 3.670 687.970 4.280 ;
        RECT 688.810 3.670 690.270 4.280 ;
        RECT 691.110 3.670 692.110 4.280 ;
        RECT 692.950 3.670 694.410 4.280 ;
        RECT 695.250 3.670 696.250 4.280 ;
        RECT 697.090 3.670 698.090 4.280 ;
        RECT 698.930 3.670 700.390 4.280 ;
        RECT 701.230 3.670 702.230 4.280 ;
        RECT 703.070 3.670 704.530 4.280 ;
        RECT 705.370 3.670 706.370 4.280 ;
        RECT 707.210 3.670 708.210 4.280 ;
        RECT 709.050 3.670 710.510 4.280 ;
        RECT 711.350 3.670 712.350 4.280 ;
        RECT 713.190 3.670 714.650 4.280 ;
        RECT 715.490 3.670 716.490 4.280 ;
        RECT 717.330 3.670 718.790 4.280 ;
        RECT 719.630 3.670 720.630 4.280 ;
        RECT 721.470 3.670 722.470 4.280 ;
        RECT 723.310 3.670 724.770 4.280 ;
        RECT 725.610 3.670 726.610 4.280 ;
        RECT 727.450 3.670 728.910 4.280 ;
        RECT 729.750 3.670 730.750 4.280 ;
        RECT 731.590 3.670 732.590 4.280 ;
        RECT 733.430 3.670 734.890 4.280 ;
        RECT 735.730 3.670 736.730 4.280 ;
        RECT 737.570 3.670 739.030 4.280 ;
        RECT 739.870 3.670 740.870 4.280 ;
        RECT 741.710 3.670 742.710 4.280 ;
        RECT 743.550 3.670 745.010 4.280 ;
        RECT 745.850 3.670 746.850 4.280 ;
        RECT 747.690 3.670 749.150 4.280 ;
        RECT 749.990 3.670 750.990 4.280 ;
        RECT 751.830 3.670 753.290 4.280 ;
        RECT 754.130 3.670 755.130 4.280 ;
        RECT 755.970 3.670 756.970 4.280 ;
        RECT 757.810 3.670 759.270 4.280 ;
        RECT 760.110 3.670 761.110 4.280 ;
        RECT 761.950 3.670 763.410 4.280 ;
        RECT 764.250 3.670 765.250 4.280 ;
        RECT 766.090 3.670 767.090 4.280 ;
        RECT 767.930 3.670 769.390 4.280 ;
        RECT 770.230 3.670 771.230 4.280 ;
        RECT 772.070 3.670 773.530 4.280 ;
        RECT 774.370 3.670 775.370 4.280 ;
        RECT 776.210 3.670 777.210 4.280 ;
        RECT 778.050 3.670 779.510 4.280 ;
        RECT 780.350 3.670 781.350 4.280 ;
        RECT 782.190 3.670 783.650 4.280 ;
        RECT 784.490 3.670 785.490 4.280 ;
        RECT 786.330 3.670 787.330 4.280 ;
        RECT 788.170 3.670 789.630 4.280 ;
        RECT 790.470 3.670 791.470 4.280 ;
        RECT 792.310 3.670 793.770 4.280 ;
        RECT 794.610 3.670 795.610 4.280 ;
        RECT 796.450 3.670 797.910 4.280 ;
        RECT 798.750 3.670 799.750 4.280 ;
        RECT 800.590 3.670 801.590 4.280 ;
        RECT 802.430 3.670 803.890 4.280 ;
        RECT 804.730 3.670 805.730 4.280 ;
        RECT 806.570 3.670 808.030 4.280 ;
        RECT 808.870 3.670 809.870 4.280 ;
        RECT 810.710 3.670 811.710 4.280 ;
        RECT 812.550 3.670 814.010 4.280 ;
        RECT 814.850 3.670 815.850 4.280 ;
        RECT 816.690 3.670 818.150 4.280 ;
        RECT 818.990 3.670 819.990 4.280 ;
        RECT 820.830 3.670 821.830 4.280 ;
        RECT 822.670 3.670 824.130 4.280 ;
        RECT 824.970 3.670 825.970 4.280 ;
        RECT 826.810 3.670 828.270 4.280 ;
        RECT 829.110 3.670 830.110 4.280 ;
        RECT 830.950 3.670 831.950 4.280 ;
        RECT 832.790 3.670 834.250 4.280 ;
        RECT 835.090 3.670 836.090 4.280 ;
        RECT 836.930 3.670 838.390 4.280 ;
        RECT 839.230 3.670 840.230 4.280 ;
        RECT 841.070 3.670 842.530 4.280 ;
        RECT 843.370 3.670 844.370 4.280 ;
        RECT 845.210 3.670 846.210 4.280 ;
        RECT 847.050 3.670 848.510 4.280 ;
        RECT 849.350 3.670 850.350 4.280 ;
        RECT 851.190 3.670 852.650 4.280 ;
        RECT 853.490 3.670 854.490 4.280 ;
        RECT 855.330 3.670 856.330 4.280 ;
        RECT 857.170 3.670 858.630 4.280 ;
        RECT 859.470 3.670 860.470 4.280 ;
        RECT 861.310 3.670 862.770 4.280 ;
        RECT 863.610 3.670 864.610 4.280 ;
        RECT 865.450 3.670 866.450 4.280 ;
        RECT 867.290 3.670 868.750 4.280 ;
        RECT 869.590 3.670 870.590 4.280 ;
        RECT 871.430 3.670 872.890 4.280 ;
        RECT 873.730 3.670 874.730 4.280 ;
        RECT 875.570 3.670 877.030 4.280 ;
        RECT 877.870 3.670 878.870 4.280 ;
        RECT 879.710 3.670 880.710 4.280 ;
        RECT 881.550 3.670 883.010 4.280 ;
        RECT 883.850 3.670 884.850 4.280 ;
        RECT 885.690 3.670 887.150 4.280 ;
        RECT 887.990 3.670 888.990 4.280 ;
        RECT 889.830 3.670 890.830 4.280 ;
        RECT 891.670 3.670 893.130 4.280 ;
        RECT 893.970 3.670 894.970 4.280 ;
        RECT 895.810 3.670 897.270 4.280 ;
        RECT 898.110 3.670 899.110 4.280 ;
        RECT 899.950 3.670 900.950 4.280 ;
        RECT 901.790 3.670 903.250 4.280 ;
        RECT 904.090 3.670 905.090 4.280 ;
        RECT 905.930 3.670 907.390 4.280 ;
        RECT 908.230 3.670 909.230 4.280 ;
        RECT 910.070 3.670 911.070 4.280 ;
        RECT 911.910 3.670 913.370 4.280 ;
        RECT 914.210 3.670 915.210 4.280 ;
        RECT 916.050 3.670 917.510 4.280 ;
        RECT 918.350 3.670 919.350 4.280 ;
        RECT 920.190 3.670 921.650 4.280 ;
        RECT 922.490 3.670 923.490 4.280 ;
        RECT 924.330 3.670 925.330 4.280 ;
        RECT 926.170 3.670 927.630 4.280 ;
        RECT 928.470 3.670 929.470 4.280 ;
        RECT 930.310 3.670 931.770 4.280 ;
        RECT 932.610 3.670 933.610 4.280 ;
        RECT 934.450 3.670 935.450 4.280 ;
        RECT 936.290 3.670 937.750 4.280 ;
        RECT 938.590 3.670 939.590 4.280 ;
        RECT 940.430 3.670 941.890 4.280 ;
        RECT 942.730 3.670 943.730 4.280 ;
        RECT 944.570 3.670 945.570 4.280 ;
        RECT 946.410 3.670 947.870 4.280 ;
        RECT 948.710 3.670 949.710 4.280 ;
        RECT 950.550 3.670 952.010 4.280 ;
        RECT 952.850 3.670 953.850 4.280 ;
        RECT 954.690 3.670 955.690 4.280 ;
        RECT 956.530 3.670 957.990 4.280 ;
        RECT 958.830 3.670 959.830 4.280 ;
        RECT 960.670 3.670 962.130 4.280 ;
        RECT 962.970 3.670 963.970 4.280 ;
        RECT 964.810 3.670 966.270 4.280 ;
        RECT 967.110 3.670 968.110 4.280 ;
        RECT 968.950 3.670 969.950 4.280 ;
        RECT 970.790 3.670 972.250 4.280 ;
        RECT 973.090 3.670 974.090 4.280 ;
        RECT 974.930 3.670 976.390 4.280 ;
        RECT 977.230 3.670 978.230 4.280 ;
        RECT 979.070 3.670 980.070 4.280 ;
        RECT 980.910 3.670 982.370 4.280 ;
        RECT 983.210 3.670 984.210 4.280 ;
        RECT 985.050 3.670 986.510 4.280 ;
        RECT 987.350 3.670 988.350 4.280 ;
        RECT 989.190 3.670 990.190 4.280 ;
        RECT 991.030 3.670 992.490 4.280 ;
        RECT 993.330 3.670 994.330 4.280 ;
        RECT 995.170 3.670 996.630 4.280 ;
        RECT 997.470 3.670 998.470 4.280 ;
      LAYER met3 ;
        RECT 0.065 10.715 944.240 987.525 ;
      LAYER met4 ;
        RECT 96.895 205.535 97.440 839.625 ;
        RECT 99.840 205.535 174.240 839.625 ;
        RECT 176.640 205.535 251.040 839.625 ;
        RECT 253.440 205.535 327.840 839.625 ;
        RECT 330.240 205.535 404.640 839.625 ;
        RECT 407.040 205.535 481.440 839.625 ;
        RECT 483.840 205.535 558.240 839.625 ;
        RECT 560.640 205.535 635.040 839.625 ;
        RECT 637.440 205.535 711.840 839.625 ;
        RECT 714.240 205.535 767.905 839.625 ;
  END
END computer
END LIBRARY

