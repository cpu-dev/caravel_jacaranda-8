magic
tech sky130A
magscale 1 2
timestamp 1634991422
<< obsli1 >>
rect 1104 2159 398820 397681
<< obsm1 >>
rect 382 1912 399634 397712
<< metal2 >>
rect 1766 399200 1822 400000
rect 5262 399200 5318 400000
rect 8758 399200 8814 400000
rect 12254 399200 12310 400000
rect 15750 399200 15806 400000
rect 19246 399200 19302 400000
rect 22742 399200 22798 400000
rect 26238 399200 26294 400000
rect 29826 399200 29882 400000
rect 33322 399200 33378 400000
rect 36818 399200 36874 400000
rect 40314 399200 40370 400000
rect 43810 399200 43866 400000
rect 47306 399200 47362 400000
rect 50802 399200 50858 400000
rect 54390 399200 54446 400000
rect 57886 399200 57942 400000
rect 61382 399200 61438 400000
rect 64878 399200 64934 400000
rect 68374 399200 68430 400000
rect 71870 399200 71926 400000
rect 75366 399200 75422 400000
rect 78954 399200 79010 400000
rect 82450 399200 82506 400000
rect 85946 399200 86002 400000
rect 89442 399200 89498 400000
rect 92938 399200 92994 400000
rect 96434 399200 96490 400000
rect 99930 399200 99986 400000
rect 103518 399200 103574 400000
rect 107014 399200 107070 400000
rect 110510 399200 110566 400000
rect 114006 399200 114062 400000
rect 117502 399200 117558 400000
rect 120998 399200 121054 400000
rect 124494 399200 124550 400000
rect 128082 399200 128138 400000
rect 131578 399200 131634 400000
rect 135074 399200 135130 400000
rect 138570 399200 138626 400000
rect 142066 399200 142122 400000
rect 145562 399200 145618 400000
rect 149058 399200 149114 400000
rect 152646 399200 152702 400000
rect 156142 399200 156198 400000
rect 159638 399200 159694 400000
rect 163134 399200 163190 400000
rect 166630 399200 166686 400000
rect 170126 399200 170182 400000
rect 173622 399200 173678 400000
rect 177210 399200 177266 400000
rect 180706 399200 180762 400000
rect 184202 399200 184258 400000
rect 187698 399200 187754 400000
rect 191194 399200 191250 400000
rect 194690 399200 194746 400000
rect 198186 399200 198242 400000
rect 201774 399200 201830 400000
rect 205270 399200 205326 400000
rect 208766 399200 208822 400000
rect 212262 399200 212318 400000
rect 215758 399200 215814 400000
rect 219254 399200 219310 400000
rect 222750 399200 222806 400000
rect 226246 399200 226302 400000
rect 229834 399200 229890 400000
rect 233330 399200 233386 400000
rect 236826 399200 236882 400000
rect 240322 399200 240378 400000
rect 243818 399200 243874 400000
rect 247314 399200 247370 400000
rect 250810 399200 250866 400000
rect 254398 399200 254454 400000
rect 257894 399200 257950 400000
rect 261390 399200 261446 400000
rect 264886 399200 264942 400000
rect 268382 399200 268438 400000
rect 271878 399200 271934 400000
rect 275374 399200 275430 400000
rect 278962 399200 279018 400000
rect 282458 399200 282514 400000
rect 285954 399200 286010 400000
rect 289450 399200 289506 400000
rect 292946 399200 293002 400000
rect 296442 399200 296498 400000
rect 299938 399200 299994 400000
rect 303526 399200 303582 400000
rect 307022 399200 307078 400000
rect 310518 399200 310574 400000
rect 314014 399200 314070 400000
rect 317510 399200 317566 400000
rect 321006 399200 321062 400000
rect 324502 399200 324558 400000
rect 328090 399200 328146 400000
rect 331586 399200 331642 400000
rect 335082 399200 335138 400000
rect 338578 399200 338634 400000
rect 342074 399200 342130 400000
rect 345570 399200 345626 400000
rect 349066 399200 349122 400000
rect 352654 399200 352710 400000
rect 356150 399200 356206 400000
rect 359646 399200 359702 400000
rect 363142 399200 363198 400000
rect 366638 399200 366694 400000
rect 370134 399200 370190 400000
rect 373630 399200 373686 400000
rect 377218 399200 377274 400000
rect 380714 399200 380770 400000
rect 384210 399200 384266 400000
rect 387706 399200 387762 400000
rect 391202 399200 391258 400000
rect 394698 399200 394754 400000
rect 398194 399200 398250 400000
rect 386 0 442 800
rect 1122 0 1178 800
rect 1950 0 2006 800
rect 2778 0 2834 800
rect 3606 0 3662 800
rect 4434 0 4490 800
rect 5170 0 5226 800
rect 5998 0 6054 800
rect 6826 0 6882 800
rect 7654 0 7710 800
rect 8482 0 8538 800
rect 9310 0 9366 800
rect 10046 0 10102 800
rect 10874 0 10930 800
rect 11702 0 11758 800
rect 12530 0 12586 800
rect 13358 0 13414 800
rect 14094 0 14150 800
rect 14922 0 14978 800
rect 15750 0 15806 800
rect 16578 0 16634 800
rect 17406 0 17462 800
rect 18234 0 18290 800
rect 18970 0 19026 800
rect 19798 0 19854 800
rect 20626 0 20682 800
rect 21454 0 21510 800
rect 22282 0 22338 800
rect 23018 0 23074 800
rect 23846 0 23902 800
rect 24674 0 24730 800
rect 25502 0 25558 800
rect 26330 0 26386 800
rect 27158 0 27214 800
rect 27894 0 27950 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30378 0 30434 800
rect 31206 0 31262 800
rect 31942 0 31998 800
rect 32770 0 32826 800
rect 33598 0 33654 800
rect 34426 0 34482 800
rect 35254 0 35310 800
rect 36082 0 36138 800
rect 36818 0 36874 800
rect 37646 0 37702 800
rect 38474 0 38530 800
rect 39302 0 39358 800
rect 40130 0 40186 800
rect 40866 0 40922 800
rect 41694 0 41750 800
rect 42522 0 42578 800
rect 43350 0 43406 800
rect 44178 0 44234 800
rect 45006 0 45062 800
rect 45742 0 45798 800
rect 46570 0 46626 800
rect 47398 0 47454 800
rect 48226 0 48282 800
rect 49054 0 49110 800
rect 49790 0 49846 800
rect 50618 0 50674 800
rect 51446 0 51502 800
rect 52274 0 52330 800
rect 53102 0 53158 800
rect 53930 0 53986 800
rect 54666 0 54722 800
rect 55494 0 55550 800
rect 56322 0 56378 800
rect 57150 0 57206 800
rect 57978 0 58034 800
rect 58806 0 58862 800
rect 59542 0 59598 800
rect 60370 0 60426 800
rect 61198 0 61254 800
rect 62026 0 62082 800
rect 62854 0 62910 800
rect 63590 0 63646 800
rect 64418 0 64474 800
rect 65246 0 65302 800
rect 66074 0 66130 800
rect 66902 0 66958 800
rect 67730 0 67786 800
rect 68466 0 68522 800
rect 69294 0 69350 800
rect 70122 0 70178 800
rect 70950 0 71006 800
rect 71778 0 71834 800
rect 72514 0 72570 800
rect 73342 0 73398 800
rect 74170 0 74226 800
rect 74998 0 75054 800
rect 75826 0 75882 800
rect 76654 0 76710 800
rect 77390 0 77446 800
rect 78218 0 78274 800
rect 79046 0 79102 800
rect 79874 0 79930 800
rect 80702 0 80758 800
rect 81438 0 81494 800
rect 82266 0 82322 800
rect 83094 0 83150 800
rect 83922 0 83978 800
rect 84750 0 84806 800
rect 85578 0 85634 800
rect 86314 0 86370 800
rect 87142 0 87198 800
rect 87970 0 88026 800
rect 88798 0 88854 800
rect 89626 0 89682 800
rect 90362 0 90418 800
rect 91190 0 91246 800
rect 92018 0 92074 800
rect 92846 0 92902 800
rect 93674 0 93730 800
rect 94502 0 94558 800
rect 95238 0 95294 800
rect 96066 0 96122 800
rect 96894 0 96950 800
rect 97722 0 97778 800
rect 98550 0 98606 800
rect 99286 0 99342 800
rect 100114 0 100170 800
rect 100942 0 100998 800
rect 101770 0 101826 800
rect 102598 0 102654 800
rect 103426 0 103482 800
rect 104162 0 104218 800
rect 104990 0 105046 800
rect 105818 0 105874 800
rect 106646 0 106702 800
rect 107474 0 107530 800
rect 108210 0 108266 800
rect 109038 0 109094 800
rect 109866 0 109922 800
rect 110694 0 110750 800
rect 111522 0 111578 800
rect 112350 0 112406 800
rect 113086 0 113142 800
rect 113914 0 113970 800
rect 114742 0 114798 800
rect 115570 0 115626 800
rect 116398 0 116454 800
rect 117226 0 117282 800
rect 117962 0 118018 800
rect 118790 0 118846 800
rect 119618 0 119674 800
rect 120446 0 120502 800
rect 121274 0 121330 800
rect 122010 0 122066 800
rect 122838 0 122894 800
rect 123666 0 123722 800
rect 124494 0 124550 800
rect 125322 0 125378 800
rect 126150 0 126206 800
rect 126886 0 126942 800
rect 127714 0 127770 800
rect 128542 0 128598 800
rect 129370 0 129426 800
rect 130198 0 130254 800
rect 130934 0 130990 800
rect 131762 0 131818 800
rect 132590 0 132646 800
rect 133418 0 133474 800
rect 134246 0 134302 800
rect 135074 0 135130 800
rect 135810 0 135866 800
rect 136638 0 136694 800
rect 137466 0 137522 800
rect 138294 0 138350 800
rect 139122 0 139178 800
rect 139858 0 139914 800
rect 140686 0 140742 800
rect 141514 0 141570 800
rect 142342 0 142398 800
rect 143170 0 143226 800
rect 143998 0 144054 800
rect 144734 0 144790 800
rect 145562 0 145618 800
rect 146390 0 146446 800
rect 147218 0 147274 800
rect 148046 0 148102 800
rect 148782 0 148838 800
rect 149610 0 149666 800
rect 150438 0 150494 800
rect 151266 0 151322 800
rect 152094 0 152150 800
rect 152922 0 152978 800
rect 153658 0 153714 800
rect 154486 0 154542 800
rect 155314 0 155370 800
rect 156142 0 156198 800
rect 156970 0 157026 800
rect 157706 0 157762 800
rect 158534 0 158590 800
rect 159362 0 159418 800
rect 160190 0 160246 800
rect 161018 0 161074 800
rect 161846 0 161902 800
rect 162582 0 162638 800
rect 163410 0 163466 800
rect 164238 0 164294 800
rect 165066 0 165122 800
rect 165894 0 165950 800
rect 166630 0 166686 800
rect 167458 0 167514 800
rect 168286 0 168342 800
rect 169114 0 169170 800
rect 169942 0 169998 800
rect 170770 0 170826 800
rect 171506 0 171562 800
rect 172334 0 172390 800
rect 173162 0 173218 800
rect 173990 0 174046 800
rect 174818 0 174874 800
rect 175646 0 175702 800
rect 176382 0 176438 800
rect 177210 0 177266 800
rect 178038 0 178094 800
rect 178866 0 178922 800
rect 179694 0 179750 800
rect 180430 0 180486 800
rect 181258 0 181314 800
rect 182086 0 182142 800
rect 182914 0 182970 800
rect 183742 0 183798 800
rect 184570 0 184626 800
rect 185306 0 185362 800
rect 186134 0 186190 800
rect 186962 0 187018 800
rect 187790 0 187846 800
rect 188618 0 188674 800
rect 189354 0 189410 800
rect 190182 0 190238 800
rect 191010 0 191066 800
rect 191838 0 191894 800
rect 192666 0 192722 800
rect 193494 0 193550 800
rect 194230 0 194286 800
rect 195058 0 195114 800
rect 195886 0 195942 800
rect 196714 0 196770 800
rect 197542 0 197598 800
rect 198278 0 198334 800
rect 199106 0 199162 800
rect 199934 0 199990 800
rect 200762 0 200818 800
rect 201590 0 201646 800
rect 202418 0 202474 800
rect 203154 0 203210 800
rect 203982 0 204038 800
rect 204810 0 204866 800
rect 205638 0 205694 800
rect 206466 0 206522 800
rect 207202 0 207258 800
rect 208030 0 208086 800
rect 208858 0 208914 800
rect 209686 0 209742 800
rect 210514 0 210570 800
rect 211342 0 211398 800
rect 212078 0 212134 800
rect 212906 0 212962 800
rect 213734 0 213790 800
rect 214562 0 214618 800
rect 215390 0 215446 800
rect 216126 0 216182 800
rect 216954 0 217010 800
rect 217782 0 217838 800
rect 218610 0 218666 800
rect 219438 0 219494 800
rect 220266 0 220322 800
rect 221002 0 221058 800
rect 221830 0 221886 800
rect 222658 0 222714 800
rect 223486 0 223542 800
rect 224314 0 224370 800
rect 225050 0 225106 800
rect 225878 0 225934 800
rect 226706 0 226762 800
rect 227534 0 227590 800
rect 228362 0 228418 800
rect 229190 0 229246 800
rect 229926 0 229982 800
rect 230754 0 230810 800
rect 231582 0 231638 800
rect 232410 0 232466 800
rect 233238 0 233294 800
rect 234066 0 234122 800
rect 234802 0 234858 800
rect 235630 0 235686 800
rect 236458 0 236514 800
rect 237286 0 237342 800
rect 238114 0 238170 800
rect 238850 0 238906 800
rect 239678 0 239734 800
rect 240506 0 240562 800
rect 241334 0 241390 800
rect 242162 0 242218 800
rect 242990 0 243046 800
rect 243726 0 243782 800
rect 244554 0 244610 800
rect 245382 0 245438 800
rect 246210 0 246266 800
rect 247038 0 247094 800
rect 247774 0 247830 800
rect 248602 0 248658 800
rect 249430 0 249486 800
rect 250258 0 250314 800
rect 251086 0 251142 800
rect 251914 0 251970 800
rect 252650 0 252706 800
rect 253478 0 253534 800
rect 254306 0 254362 800
rect 255134 0 255190 800
rect 255962 0 256018 800
rect 256698 0 256754 800
rect 257526 0 257582 800
rect 258354 0 258410 800
rect 259182 0 259238 800
rect 260010 0 260066 800
rect 260838 0 260894 800
rect 261574 0 261630 800
rect 262402 0 262458 800
rect 263230 0 263286 800
rect 264058 0 264114 800
rect 264886 0 264942 800
rect 265622 0 265678 800
rect 266450 0 266506 800
rect 267278 0 267334 800
rect 268106 0 268162 800
rect 268934 0 268990 800
rect 269762 0 269818 800
rect 270498 0 270554 800
rect 271326 0 271382 800
rect 272154 0 272210 800
rect 272982 0 273038 800
rect 273810 0 273866 800
rect 274546 0 274602 800
rect 275374 0 275430 800
rect 276202 0 276258 800
rect 277030 0 277086 800
rect 277858 0 277914 800
rect 278686 0 278742 800
rect 279422 0 279478 800
rect 280250 0 280306 800
rect 281078 0 281134 800
rect 281906 0 281962 800
rect 282734 0 282790 800
rect 283470 0 283526 800
rect 284298 0 284354 800
rect 285126 0 285182 800
rect 285954 0 286010 800
rect 286782 0 286838 800
rect 287610 0 287666 800
rect 288346 0 288402 800
rect 289174 0 289230 800
rect 290002 0 290058 800
rect 290830 0 290886 800
rect 291658 0 291714 800
rect 292486 0 292542 800
rect 293222 0 293278 800
rect 294050 0 294106 800
rect 294878 0 294934 800
rect 295706 0 295762 800
rect 296534 0 296590 800
rect 297270 0 297326 800
rect 298098 0 298154 800
rect 298926 0 298982 800
rect 299754 0 299810 800
rect 300582 0 300638 800
rect 301410 0 301466 800
rect 302146 0 302202 800
rect 302974 0 303030 800
rect 303802 0 303858 800
rect 304630 0 304686 800
rect 305458 0 305514 800
rect 306194 0 306250 800
rect 307022 0 307078 800
rect 307850 0 307906 800
rect 308678 0 308734 800
rect 309506 0 309562 800
rect 310334 0 310390 800
rect 311070 0 311126 800
rect 311898 0 311954 800
rect 312726 0 312782 800
rect 313554 0 313610 800
rect 314382 0 314438 800
rect 315118 0 315174 800
rect 315946 0 316002 800
rect 316774 0 316830 800
rect 317602 0 317658 800
rect 318430 0 318486 800
rect 319258 0 319314 800
rect 319994 0 320050 800
rect 320822 0 320878 800
rect 321650 0 321706 800
rect 322478 0 322534 800
rect 323306 0 323362 800
rect 324042 0 324098 800
rect 324870 0 324926 800
rect 325698 0 325754 800
rect 326526 0 326582 800
rect 327354 0 327410 800
rect 328182 0 328238 800
rect 328918 0 328974 800
rect 329746 0 329802 800
rect 330574 0 330630 800
rect 331402 0 331458 800
rect 332230 0 332286 800
rect 332966 0 333022 800
rect 333794 0 333850 800
rect 334622 0 334678 800
rect 335450 0 335506 800
rect 336278 0 336334 800
rect 337106 0 337162 800
rect 337842 0 337898 800
rect 338670 0 338726 800
rect 339498 0 339554 800
rect 340326 0 340382 800
rect 341154 0 341210 800
rect 341890 0 341946 800
rect 342718 0 342774 800
rect 343546 0 343602 800
rect 344374 0 344430 800
rect 345202 0 345258 800
rect 346030 0 346086 800
rect 346766 0 346822 800
rect 347594 0 347650 800
rect 348422 0 348478 800
rect 349250 0 349306 800
rect 350078 0 350134 800
rect 350906 0 350962 800
rect 351642 0 351698 800
rect 352470 0 352526 800
rect 353298 0 353354 800
rect 354126 0 354182 800
rect 354954 0 355010 800
rect 355690 0 355746 800
rect 356518 0 356574 800
rect 357346 0 357402 800
rect 358174 0 358230 800
rect 359002 0 359058 800
rect 359830 0 359886 800
rect 360566 0 360622 800
rect 361394 0 361450 800
rect 362222 0 362278 800
rect 363050 0 363106 800
rect 363878 0 363934 800
rect 364614 0 364670 800
rect 365442 0 365498 800
rect 366270 0 366326 800
rect 367098 0 367154 800
rect 367926 0 367982 800
rect 368754 0 368810 800
rect 369490 0 369546 800
rect 370318 0 370374 800
rect 371146 0 371202 800
rect 371974 0 372030 800
rect 372802 0 372858 800
rect 373538 0 373594 800
rect 374366 0 374422 800
rect 375194 0 375250 800
rect 376022 0 376078 800
rect 376850 0 376906 800
rect 377678 0 377734 800
rect 378414 0 378470 800
rect 379242 0 379298 800
rect 380070 0 380126 800
rect 380898 0 380954 800
rect 381726 0 381782 800
rect 382462 0 382518 800
rect 383290 0 383346 800
rect 384118 0 384174 800
rect 384946 0 385002 800
rect 385774 0 385830 800
rect 386602 0 386658 800
rect 387338 0 387394 800
rect 388166 0 388222 800
rect 388994 0 389050 800
rect 389822 0 389878 800
rect 390650 0 390706 800
rect 391386 0 391442 800
rect 392214 0 392270 800
rect 393042 0 393098 800
rect 393870 0 393926 800
rect 394698 0 394754 800
rect 395526 0 395582 800
rect 396262 0 396318 800
rect 397090 0 397146 800
rect 397918 0 397974 800
rect 398746 0 398802 800
rect 399574 0 399630 800
<< obsm2 >>
rect 388 399144 1710 399242
rect 1878 399144 5206 399242
rect 5374 399144 8702 399242
rect 8870 399144 12198 399242
rect 12366 399144 15694 399242
rect 15862 399144 19190 399242
rect 19358 399144 22686 399242
rect 22854 399144 26182 399242
rect 26350 399144 29770 399242
rect 29938 399144 33266 399242
rect 33434 399144 36762 399242
rect 36930 399144 40258 399242
rect 40426 399144 43754 399242
rect 43922 399144 47250 399242
rect 47418 399144 50746 399242
rect 50914 399144 54334 399242
rect 54502 399144 57830 399242
rect 57998 399144 61326 399242
rect 61494 399144 64822 399242
rect 64990 399144 68318 399242
rect 68486 399144 71814 399242
rect 71982 399144 75310 399242
rect 75478 399144 78898 399242
rect 79066 399144 82394 399242
rect 82562 399144 85890 399242
rect 86058 399144 89386 399242
rect 89554 399144 92882 399242
rect 93050 399144 96378 399242
rect 96546 399144 99874 399242
rect 100042 399144 103462 399242
rect 103630 399144 106958 399242
rect 107126 399144 110454 399242
rect 110622 399144 113950 399242
rect 114118 399144 117446 399242
rect 117614 399144 120942 399242
rect 121110 399144 124438 399242
rect 124606 399144 128026 399242
rect 128194 399144 131522 399242
rect 131690 399144 135018 399242
rect 135186 399144 138514 399242
rect 138682 399144 142010 399242
rect 142178 399144 145506 399242
rect 145674 399144 149002 399242
rect 149170 399144 152590 399242
rect 152758 399144 156086 399242
rect 156254 399144 159582 399242
rect 159750 399144 163078 399242
rect 163246 399144 166574 399242
rect 166742 399144 170070 399242
rect 170238 399144 173566 399242
rect 173734 399144 177154 399242
rect 177322 399144 180650 399242
rect 180818 399144 184146 399242
rect 184314 399144 187642 399242
rect 187810 399144 191138 399242
rect 191306 399144 194634 399242
rect 194802 399144 198130 399242
rect 198298 399144 201718 399242
rect 201886 399144 205214 399242
rect 205382 399144 208710 399242
rect 208878 399144 212206 399242
rect 212374 399144 215702 399242
rect 215870 399144 219198 399242
rect 219366 399144 222694 399242
rect 222862 399144 226190 399242
rect 226358 399144 229778 399242
rect 229946 399144 233274 399242
rect 233442 399144 236770 399242
rect 236938 399144 240266 399242
rect 240434 399144 243762 399242
rect 243930 399144 247258 399242
rect 247426 399144 250754 399242
rect 250922 399144 254342 399242
rect 254510 399144 257838 399242
rect 258006 399144 261334 399242
rect 261502 399144 264830 399242
rect 264998 399144 268326 399242
rect 268494 399144 271822 399242
rect 271990 399144 275318 399242
rect 275486 399144 278906 399242
rect 279074 399144 282402 399242
rect 282570 399144 285898 399242
rect 286066 399144 289394 399242
rect 289562 399144 292890 399242
rect 293058 399144 296386 399242
rect 296554 399144 299882 399242
rect 300050 399144 303470 399242
rect 303638 399144 306966 399242
rect 307134 399144 310462 399242
rect 310630 399144 313958 399242
rect 314126 399144 317454 399242
rect 317622 399144 320950 399242
rect 321118 399144 324446 399242
rect 324614 399144 328034 399242
rect 328202 399144 331530 399242
rect 331698 399144 335026 399242
rect 335194 399144 338522 399242
rect 338690 399144 342018 399242
rect 342186 399144 345514 399242
rect 345682 399144 349010 399242
rect 349178 399144 352598 399242
rect 352766 399144 356094 399242
rect 356262 399144 359590 399242
rect 359758 399144 363086 399242
rect 363254 399144 366582 399242
rect 366750 399144 370078 399242
rect 370246 399144 373574 399242
rect 373742 399144 377162 399242
rect 377330 399144 380658 399242
rect 380826 399144 384154 399242
rect 384322 399144 387650 399242
rect 387818 399144 391146 399242
rect 391314 399144 394642 399242
rect 394810 399144 398138 399242
rect 398306 399144 399628 399242
rect 388 856 399628 399144
rect 498 734 1066 856
rect 1234 734 1894 856
rect 2062 734 2722 856
rect 2890 734 3550 856
rect 3718 734 4378 856
rect 4546 734 5114 856
rect 5282 734 5942 856
rect 6110 734 6770 856
rect 6938 734 7598 856
rect 7766 734 8426 856
rect 8594 734 9254 856
rect 9422 734 9990 856
rect 10158 734 10818 856
rect 10986 734 11646 856
rect 11814 734 12474 856
rect 12642 734 13302 856
rect 13470 734 14038 856
rect 14206 734 14866 856
rect 15034 734 15694 856
rect 15862 734 16522 856
rect 16690 734 17350 856
rect 17518 734 18178 856
rect 18346 734 18914 856
rect 19082 734 19742 856
rect 19910 734 20570 856
rect 20738 734 21398 856
rect 21566 734 22226 856
rect 22394 734 22962 856
rect 23130 734 23790 856
rect 23958 734 24618 856
rect 24786 734 25446 856
rect 25614 734 26274 856
rect 26442 734 27102 856
rect 27270 734 27838 856
rect 28006 734 28666 856
rect 28834 734 29494 856
rect 29662 734 30322 856
rect 30490 734 31150 856
rect 31318 734 31886 856
rect 32054 734 32714 856
rect 32882 734 33542 856
rect 33710 734 34370 856
rect 34538 734 35198 856
rect 35366 734 36026 856
rect 36194 734 36762 856
rect 36930 734 37590 856
rect 37758 734 38418 856
rect 38586 734 39246 856
rect 39414 734 40074 856
rect 40242 734 40810 856
rect 40978 734 41638 856
rect 41806 734 42466 856
rect 42634 734 43294 856
rect 43462 734 44122 856
rect 44290 734 44950 856
rect 45118 734 45686 856
rect 45854 734 46514 856
rect 46682 734 47342 856
rect 47510 734 48170 856
rect 48338 734 48998 856
rect 49166 734 49734 856
rect 49902 734 50562 856
rect 50730 734 51390 856
rect 51558 734 52218 856
rect 52386 734 53046 856
rect 53214 734 53874 856
rect 54042 734 54610 856
rect 54778 734 55438 856
rect 55606 734 56266 856
rect 56434 734 57094 856
rect 57262 734 57922 856
rect 58090 734 58750 856
rect 58918 734 59486 856
rect 59654 734 60314 856
rect 60482 734 61142 856
rect 61310 734 61970 856
rect 62138 734 62798 856
rect 62966 734 63534 856
rect 63702 734 64362 856
rect 64530 734 65190 856
rect 65358 734 66018 856
rect 66186 734 66846 856
rect 67014 734 67674 856
rect 67842 734 68410 856
rect 68578 734 69238 856
rect 69406 734 70066 856
rect 70234 734 70894 856
rect 71062 734 71722 856
rect 71890 734 72458 856
rect 72626 734 73286 856
rect 73454 734 74114 856
rect 74282 734 74942 856
rect 75110 734 75770 856
rect 75938 734 76598 856
rect 76766 734 77334 856
rect 77502 734 78162 856
rect 78330 734 78990 856
rect 79158 734 79818 856
rect 79986 734 80646 856
rect 80814 734 81382 856
rect 81550 734 82210 856
rect 82378 734 83038 856
rect 83206 734 83866 856
rect 84034 734 84694 856
rect 84862 734 85522 856
rect 85690 734 86258 856
rect 86426 734 87086 856
rect 87254 734 87914 856
rect 88082 734 88742 856
rect 88910 734 89570 856
rect 89738 734 90306 856
rect 90474 734 91134 856
rect 91302 734 91962 856
rect 92130 734 92790 856
rect 92958 734 93618 856
rect 93786 734 94446 856
rect 94614 734 95182 856
rect 95350 734 96010 856
rect 96178 734 96838 856
rect 97006 734 97666 856
rect 97834 734 98494 856
rect 98662 734 99230 856
rect 99398 734 100058 856
rect 100226 734 100886 856
rect 101054 734 101714 856
rect 101882 734 102542 856
rect 102710 734 103370 856
rect 103538 734 104106 856
rect 104274 734 104934 856
rect 105102 734 105762 856
rect 105930 734 106590 856
rect 106758 734 107418 856
rect 107586 734 108154 856
rect 108322 734 108982 856
rect 109150 734 109810 856
rect 109978 734 110638 856
rect 110806 734 111466 856
rect 111634 734 112294 856
rect 112462 734 113030 856
rect 113198 734 113858 856
rect 114026 734 114686 856
rect 114854 734 115514 856
rect 115682 734 116342 856
rect 116510 734 117170 856
rect 117338 734 117906 856
rect 118074 734 118734 856
rect 118902 734 119562 856
rect 119730 734 120390 856
rect 120558 734 121218 856
rect 121386 734 121954 856
rect 122122 734 122782 856
rect 122950 734 123610 856
rect 123778 734 124438 856
rect 124606 734 125266 856
rect 125434 734 126094 856
rect 126262 734 126830 856
rect 126998 734 127658 856
rect 127826 734 128486 856
rect 128654 734 129314 856
rect 129482 734 130142 856
rect 130310 734 130878 856
rect 131046 734 131706 856
rect 131874 734 132534 856
rect 132702 734 133362 856
rect 133530 734 134190 856
rect 134358 734 135018 856
rect 135186 734 135754 856
rect 135922 734 136582 856
rect 136750 734 137410 856
rect 137578 734 138238 856
rect 138406 734 139066 856
rect 139234 734 139802 856
rect 139970 734 140630 856
rect 140798 734 141458 856
rect 141626 734 142286 856
rect 142454 734 143114 856
rect 143282 734 143942 856
rect 144110 734 144678 856
rect 144846 734 145506 856
rect 145674 734 146334 856
rect 146502 734 147162 856
rect 147330 734 147990 856
rect 148158 734 148726 856
rect 148894 734 149554 856
rect 149722 734 150382 856
rect 150550 734 151210 856
rect 151378 734 152038 856
rect 152206 734 152866 856
rect 153034 734 153602 856
rect 153770 734 154430 856
rect 154598 734 155258 856
rect 155426 734 156086 856
rect 156254 734 156914 856
rect 157082 734 157650 856
rect 157818 734 158478 856
rect 158646 734 159306 856
rect 159474 734 160134 856
rect 160302 734 160962 856
rect 161130 734 161790 856
rect 161958 734 162526 856
rect 162694 734 163354 856
rect 163522 734 164182 856
rect 164350 734 165010 856
rect 165178 734 165838 856
rect 166006 734 166574 856
rect 166742 734 167402 856
rect 167570 734 168230 856
rect 168398 734 169058 856
rect 169226 734 169886 856
rect 170054 734 170714 856
rect 170882 734 171450 856
rect 171618 734 172278 856
rect 172446 734 173106 856
rect 173274 734 173934 856
rect 174102 734 174762 856
rect 174930 734 175590 856
rect 175758 734 176326 856
rect 176494 734 177154 856
rect 177322 734 177982 856
rect 178150 734 178810 856
rect 178978 734 179638 856
rect 179806 734 180374 856
rect 180542 734 181202 856
rect 181370 734 182030 856
rect 182198 734 182858 856
rect 183026 734 183686 856
rect 183854 734 184514 856
rect 184682 734 185250 856
rect 185418 734 186078 856
rect 186246 734 186906 856
rect 187074 734 187734 856
rect 187902 734 188562 856
rect 188730 734 189298 856
rect 189466 734 190126 856
rect 190294 734 190954 856
rect 191122 734 191782 856
rect 191950 734 192610 856
rect 192778 734 193438 856
rect 193606 734 194174 856
rect 194342 734 195002 856
rect 195170 734 195830 856
rect 195998 734 196658 856
rect 196826 734 197486 856
rect 197654 734 198222 856
rect 198390 734 199050 856
rect 199218 734 199878 856
rect 200046 734 200706 856
rect 200874 734 201534 856
rect 201702 734 202362 856
rect 202530 734 203098 856
rect 203266 734 203926 856
rect 204094 734 204754 856
rect 204922 734 205582 856
rect 205750 734 206410 856
rect 206578 734 207146 856
rect 207314 734 207974 856
rect 208142 734 208802 856
rect 208970 734 209630 856
rect 209798 734 210458 856
rect 210626 734 211286 856
rect 211454 734 212022 856
rect 212190 734 212850 856
rect 213018 734 213678 856
rect 213846 734 214506 856
rect 214674 734 215334 856
rect 215502 734 216070 856
rect 216238 734 216898 856
rect 217066 734 217726 856
rect 217894 734 218554 856
rect 218722 734 219382 856
rect 219550 734 220210 856
rect 220378 734 220946 856
rect 221114 734 221774 856
rect 221942 734 222602 856
rect 222770 734 223430 856
rect 223598 734 224258 856
rect 224426 734 224994 856
rect 225162 734 225822 856
rect 225990 734 226650 856
rect 226818 734 227478 856
rect 227646 734 228306 856
rect 228474 734 229134 856
rect 229302 734 229870 856
rect 230038 734 230698 856
rect 230866 734 231526 856
rect 231694 734 232354 856
rect 232522 734 233182 856
rect 233350 734 234010 856
rect 234178 734 234746 856
rect 234914 734 235574 856
rect 235742 734 236402 856
rect 236570 734 237230 856
rect 237398 734 238058 856
rect 238226 734 238794 856
rect 238962 734 239622 856
rect 239790 734 240450 856
rect 240618 734 241278 856
rect 241446 734 242106 856
rect 242274 734 242934 856
rect 243102 734 243670 856
rect 243838 734 244498 856
rect 244666 734 245326 856
rect 245494 734 246154 856
rect 246322 734 246982 856
rect 247150 734 247718 856
rect 247886 734 248546 856
rect 248714 734 249374 856
rect 249542 734 250202 856
rect 250370 734 251030 856
rect 251198 734 251858 856
rect 252026 734 252594 856
rect 252762 734 253422 856
rect 253590 734 254250 856
rect 254418 734 255078 856
rect 255246 734 255906 856
rect 256074 734 256642 856
rect 256810 734 257470 856
rect 257638 734 258298 856
rect 258466 734 259126 856
rect 259294 734 259954 856
rect 260122 734 260782 856
rect 260950 734 261518 856
rect 261686 734 262346 856
rect 262514 734 263174 856
rect 263342 734 264002 856
rect 264170 734 264830 856
rect 264998 734 265566 856
rect 265734 734 266394 856
rect 266562 734 267222 856
rect 267390 734 268050 856
rect 268218 734 268878 856
rect 269046 734 269706 856
rect 269874 734 270442 856
rect 270610 734 271270 856
rect 271438 734 272098 856
rect 272266 734 272926 856
rect 273094 734 273754 856
rect 273922 734 274490 856
rect 274658 734 275318 856
rect 275486 734 276146 856
rect 276314 734 276974 856
rect 277142 734 277802 856
rect 277970 734 278630 856
rect 278798 734 279366 856
rect 279534 734 280194 856
rect 280362 734 281022 856
rect 281190 734 281850 856
rect 282018 734 282678 856
rect 282846 734 283414 856
rect 283582 734 284242 856
rect 284410 734 285070 856
rect 285238 734 285898 856
rect 286066 734 286726 856
rect 286894 734 287554 856
rect 287722 734 288290 856
rect 288458 734 289118 856
rect 289286 734 289946 856
rect 290114 734 290774 856
rect 290942 734 291602 856
rect 291770 734 292430 856
rect 292598 734 293166 856
rect 293334 734 293994 856
rect 294162 734 294822 856
rect 294990 734 295650 856
rect 295818 734 296478 856
rect 296646 734 297214 856
rect 297382 734 298042 856
rect 298210 734 298870 856
rect 299038 734 299698 856
rect 299866 734 300526 856
rect 300694 734 301354 856
rect 301522 734 302090 856
rect 302258 734 302918 856
rect 303086 734 303746 856
rect 303914 734 304574 856
rect 304742 734 305402 856
rect 305570 734 306138 856
rect 306306 734 306966 856
rect 307134 734 307794 856
rect 307962 734 308622 856
rect 308790 734 309450 856
rect 309618 734 310278 856
rect 310446 734 311014 856
rect 311182 734 311842 856
rect 312010 734 312670 856
rect 312838 734 313498 856
rect 313666 734 314326 856
rect 314494 734 315062 856
rect 315230 734 315890 856
rect 316058 734 316718 856
rect 316886 734 317546 856
rect 317714 734 318374 856
rect 318542 734 319202 856
rect 319370 734 319938 856
rect 320106 734 320766 856
rect 320934 734 321594 856
rect 321762 734 322422 856
rect 322590 734 323250 856
rect 323418 734 323986 856
rect 324154 734 324814 856
rect 324982 734 325642 856
rect 325810 734 326470 856
rect 326638 734 327298 856
rect 327466 734 328126 856
rect 328294 734 328862 856
rect 329030 734 329690 856
rect 329858 734 330518 856
rect 330686 734 331346 856
rect 331514 734 332174 856
rect 332342 734 332910 856
rect 333078 734 333738 856
rect 333906 734 334566 856
rect 334734 734 335394 856
rect 335562 734 336222 856
rect 336390 734 337050 856
rect 337218 734 337786 856
rect 337954 734 338614 856
rect 338782 734 339442 856
rect 339610 734 340270 856
rect 340438 734 341098 856
rect 341266 734 341834 856
rect 342002 734 342662 856
rect 342830 734 343490 856
rect 343658 734 344318 856
rect 344486 734 345146 856
rect 345314 734 345974 856
rect 346142 734 346710 856
rect 346878 734 347538 856
rect 347706 734 348366 856
rect 348534 734 349194 856
rect 349362 734 350022 856
rect 350190 734 350850 856
rect 351018 734 351586 856
rect 351754 734 352414 856
rect 352582 734 353242 856
rect 353410 734 354070 856
rect 354238 734 354898 856
rect 355066 734 355634 856
rect 355802 734 356462 856
rect 356630 734 357290 856
rect 357458 734 358118 856
rect 358286 734 358946 856
rect 359114 734 359774 856
rect 359942 734 360510 856
rect 360678 734 361338 856
rect 361506 734 362166 856
rect 362334 734 362994 856
rect 363162 734 363822 856
rect 363990 734 364558 856
rect 364726 734 365386 856
rect 365554 734 366214 856
rect 366382 734 367042 856
rect 367210 734 367870 856
rect 368038 734 368698 856
rect 368866 734 369434 856
rect 369602 734 370262 856
rect 370430 734 371090 856
rect 371258 734 371918 856
rect 372086 734 372746 856
rect 372914 734 373482 856
rect 373650 734 374310 856
rect 374478 734 375138 856
rect 375306 734 375966 856
rect 376134 734 376794 856
rect 376962 734 377622 856
rect 377790 734 378358 856
rect 378526 734 379186 856
rect 379354 734 380014 856
rect 380182 734 380842 856
rect 381010 734 381670 856
rect 381838 734 382406 856
rect 382574 734 383234 856
rect 383402 734 384062 856
rect 384230 734 384890 856
rect 385058 734 385718 856
rect 385886 734 386546 856
rect 386714 734 387282 856
rect 387450 734 388110 856
rect 388278 734 388938 856
rect 389106 734 389766 856
rect 389934 734 390594 856
rect 390762 734 391330 856
rect 391498 734 392158 856
rect 392326 734 392986 856
rect 393154 734 393814 856
rect 393982 734 394642 856
rect 394810 734 395470 856
rect 395638 734 396206 856
rect 396374 734 397034 856
rect 397202 734 397862 856
rect 398030 734 398690 856
rect 398858 734 399518 856
<< obsm3 >>
rect 4208 2143 388528 397697
<< metal4 >>
rect 4208 2128 4528 397712
rect 19568 2128 19888 397712
rect 34928 2128 35248 397712
rect 50288 2128 50608 397712
rect 65648 2128 65968 397712
rect 81008 2128 81328 397712
rect 96368 2128 96688 397712
rect 111728 2128 112048 397712
rect 127088 2128 127408 397712
rect 142448 2128 142768 397712
rect 157808 2128 158128 397712
rect 173168 2128 173488 397712
rect 188528 2128 188848 397712
rect 203888 2128 204208 397712
rect 219248 2128 219568 397712
rect 234608 2128 234928 397712
rect 249968 2128 250288 397712
rect 265328 2128 265648 397712
rect 280688 2128 281008 397712
rect 296048 2128 296368 397712
rect 311408 2128 311728 397712
rect 326768 2128 327088 397712
rect 342128 2128 342448 397712
rect 357488 2128 357808 397712
rect 372848 2128 373168 397712
rect 388208 2128 388528 397712
<< obsm4 >>
rect 50843 40019 65568 169829
rect 66048 40019 80928 169829
rect 81408 40019 96288 169829
rect 96768 40019 111648 169829
rect 112128 40019 127008 169829
rect 127488 40019 142368 169829
rect 142848 40019 157728 169829
rect 158208 40019 173088 169829
rect 173568 40019 187621 169829
<< labels >>
rlabel metal2 s 1766 399200 1822 400000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 107014 399200 107070 400000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 117502 399200 117558 400000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 128082 399200 128138 400000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 138570 399200 138626 400000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 149058 399200 149114 400000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 159638 399200 159694 400000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 170126 399200 170182 400000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 180706 399200 180762 400000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 191194 399200 191250 400000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 201774 399200 201830 400000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 12254 399200 12310 400000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 212262 399200 212318 400000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 222750 399200 222806 400000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 233330 399200 233386 400000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 243818 399200 243874 400000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 254398 399200 254454 400000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 264886 399200 264942 400000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 275374 399200 275430 400000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 285954 399200 286010 400000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 296442 399200 296498 400000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 307022 399200 307078 400000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 22742 399200 22798 400000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 317510 399200 317566 400000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 328090 399200 328146 400000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 338578 399200 338634 400000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 349066 399200 349122 400000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 359646 399200 359702 400000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 370134 399200 370190 400000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 380714 399200 380770 400000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 391202 399200 391258 400000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 33322 399200 33378 400000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 43810 399200 43866 400000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 54390 399200 54446 400000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 64878 399200 64934 400000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 75366 399200 75422 400000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 85946 399200 86002 400000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 96434 399200 96490 400000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5262 399200 5318 400000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 110510 399200 110566 400000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 120998 399200 121054 400000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 131578 399200 131634 400000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 142066 399200 142122 400000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 152646 399200 152702 400000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 163134 399200 163190 400000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 173622 399200 173678 400000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 184202 399200 184258 400000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 194690 399200 194746 400000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 205270 399200 205326 400000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 15750 399200 15806 400000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 215758 399200 215814 400000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 226246 399200 226302 400000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 236826 399200 236882 400000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 247314 399200 247370 400000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 257894 399200 257950 400000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 268382 399200 268438 400000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 278962 399200 279018 400000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 289450 399200 289506 400000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 299938 399200 299994 400000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 310518 399200 310574 400000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 26238 399200 26294 400000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 321006 399200 321062 400000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 331586 399200 331642 400000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 342074 399200 342130 400000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 352654 399200 352710 400000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 363142 399200 363198 400000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 373630 399200 373686 400000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 384210 399200 384266 400000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 394698 399200 394754 400000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 36818 399200 36874 400000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 47306 399200 47362 400000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 57886 399200 57942 400000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 68374 399200 68430 400000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 78954 399200 79010 400000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 89442 399200 89498 400000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 99930 399200 99986 400000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 8758 399200 8814 400000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 114006 399200 114062 400000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 124494 399200 124550 400000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 135074 399200 135130 400000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 145562 399200 145618 400000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 156142 399200 156198 400000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 166630 399200 166686 400000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 177210 399200 177266 400000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 187698 399200 187754 400000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 198186 399200 198242 400000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 208766 399200 208822 400000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 19246 399200 19302 400000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 219254 399200 219310 400000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 229834 399200 229890 400000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 240322 399200 240378 400000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 250810 399200 250866 400000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 261390 399200 261446 400000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 271878 399200 271934 400000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 282458 399200 282514 400000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 292946 399200 293002 400000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 303526 399200 303582 400000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 314014 399200 314070 400000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 29826 399200 29882 400000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 324502 399200 324558 400000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 335082 399200 335138 400000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 345570 399200 345626 400000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 356150 399200 356206 400000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 366638 399200 366694 400000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 377218 399200 377274 400000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 387706 399200 387762 400000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 398194 399200 398250 400000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 40314 399200 40370 400000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 50802 399200 50858 400000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 61382 399200 61438 400000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 71870 399200 71926 400000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 82450 399200 82506 400000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 92938 399200 92994 400000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 103518 399200 103574 400000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 397918 0 397974 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 398746 0 398802 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 399574 0 399630 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 329746 0 329802 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 332230 0 332286 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 334622 0 334678 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 337106 0 337162 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 339498 0 339554 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 341890 0 341946 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 344374 0 344430 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 346766 0 346822 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 349250 0 349306 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 351642 0 351698 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 354126 0 354182 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 356518 0 356574 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 359002 0 359058 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 361394 0 361450 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 363878 0 363934 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 366270 0 366326 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 368754 0 368810 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 371146 0 371202 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 373538 0 373594 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 376022 0 376078 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 378414 0 378470 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 380898 0 380954 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 383290 0 383346 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 385774 0 385830 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 388166 0 388222 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 390650 0 390706 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 393042 0 393098 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 395526 0 395582 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 176382 0 176438 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 181258 0 181314 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 198278 0 198334 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 200762 0 200818 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 203154 0 203210 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 205638 0 205694 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 217782 0 217838 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 220266 0 220322 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 227534 0 227590 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 232410 0 232466 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 237286 0 237342 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 242162 0 242218 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 244554 0 244610 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 247038 0 247094 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 249430 0 249486 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 251914 0 251970 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 254306 0 254362 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 256698 0 256754 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 259182 0 259238 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 261574 0 261630 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 264058 0 264114 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 266450 0 266506 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 268934 0 268990 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 271326 0 271382 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 273810 0 273866 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 276202 0 276258 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 278686 0 278742 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 283470 0 283526 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 285954 0 286010 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 288346 0 288402 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 290830 0 290886 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 293222 0 293278 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 295706 0 295762 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 298098 0 298154 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 300582 0 300638 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 302974 0 303030 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 305458 0 305514 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 307850 0 307906 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 310334 0 310390 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 312726 0 312782 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 315118 0 315174 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 317602 0 317658 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 319994 0 320050 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 322478 0 322534 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 324870 0 324926 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 327354 0 327410 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 330574 0 330630 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 332966 0 333022 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 335450 0 335506 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 337842 0 337898 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 340326 0 340382 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 342718 0 342774 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 345202 0 345258 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 347594 0 347650 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 350078 0 350134 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 352470 0 352526 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 354954 0 355010 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 357346 0 357402 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 359830 0 359886 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 362222 0 362278 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 364614 0 364670 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 367098 0 367154 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 369490 0 369546 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 371974 0 372030 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 374366 0 374422 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 376850 0 376906 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 379242 0 379298 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 381726 0 381782 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 384118 0 384174 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 386602 0 386658 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 388994 0 389050 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 391386 0 391442 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 393870 0 393926 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 396262 0 396318 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 130934 0 130990 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 140686 0 140742 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 143170 0 143226 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 148046 0 148102 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 157706 0 157762 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 160190 0 160246 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 162582 0 162638 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 165066 0 165122 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 172334 0 172390 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 182086 0 182142 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 184570 0 184626 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 186962 0 187018 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 189354 0 189410 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 191838 0 191894 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 194230 0 194286 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 199106 0 199162 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 201590 0 201646 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 203982 0 204038 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 206466 0 206522 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 208858 0 208914 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 211342 0 211398 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 213734 0 213790 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 216126 0 216182 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 218610 0 218666 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 221002 0 221058 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 223486 0 223542 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 225878 0 225934 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 228362 0 228418 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 230754 0 230810 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 233238 0 233294 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 235630 0 235686 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 238114 0 238170 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 240506 0 240562 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 242990 0 243046 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 245382 0 245438 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 247774 0 247830 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 250258 0 250314 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 252650 0 252706 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 255134 0 255190 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 257526 0 257582 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 260010 0 260066 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 262402 0 262458 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 264886 0 264942 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 267278 0 267334 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 269762 0 269818 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 272154 0 272210 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 274546 0 274602 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 277030 0 277086 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 279422 0 279478 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 281906 0 281962 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 284298 0 284354 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 286782 0 286838 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 289174 0 289230 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 291658 0 291714 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 294050 0 294106 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 296534 0 296590 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 298926 0 298982 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 301410 0 301466 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 303802 0 303858 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 306194 0 306250 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 308678 0 308734 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 311070 0 311126 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 313554 0 313610 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 315946 0 316002 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 318430 0 318486 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 320822 0 320878 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 323306 0 323362 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 325698 0 325754 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 328182 0 328238 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 87970 0 88026 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 331402 0 331458 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 333794 0 333850 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 336278 0 336334 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 338670 0 338726 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 341154 0 341210 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 343546 0 343602 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 346030 0 346086 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 348422 0 348478 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 350906 0 350962 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 353298 0 353354 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 355690 0 355746 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 358174 0 358230 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 360566 0 360622 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 363050 0 363106 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 365442 0 365498 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 367926 0 367982 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 370318 0 370374 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 372802 0 372858 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 375194 0 375250 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 377678 0 377734 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 380070 0 380126 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 382462 0 382518 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 384946 0 385002 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 387338 0 387394 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 389822 0 389878 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 392214 0 392270 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 394698 0 394754 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 397090 0 397146 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 175646 0 175702 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 180430 0 180486 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 185306 0 185362 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 190182 0 190238 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 192666 0 192722 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 202418 0 202474 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 209686 0 209742 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 212078 0 212134 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 214562 0 214618 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 216954 0 217010 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 219438 0 219494 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 221830 0 221886 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 224314 0 224370 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 226706 0 226762 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 229190 0 229246 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 234066 0 234122 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 236458 0 236514 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 241334 0 241390 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 243726 0 243782 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 246210 0 246266 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 251086 0 251142 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 253478 0 253534 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 258354 0 258410 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 260838 0 260894 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 263230 0 263286 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 265622 0 265678 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 268106 0 268162 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 270498 0 270554 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 272982 0 273038 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 275374 0 275430 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 277858 0 277914 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 280250 0 280306 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 282734 0 282790 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 285126 0 285182 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 287610 0 287666 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 290002 0 290058 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 292486 0 292542 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 294878 0 294934 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 297270 0 297326 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 299754 0 299810 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 302146 0 302202 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 304630 0 304686 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 307022 0 307078 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 309506 0 309562 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 311898 0 311954 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 314382 0 314438 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 316774 0 316830 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 319258 0 319314 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 321650 0 321706 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 324042 0 324098 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 326526 0 326582 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 328918 0 328974 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 397712 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 397712 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 397712 6 vssd1
port 503 nsew ground input
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 400000 400000
string LEFview TRUE
string GDS_FILE /project/openlane/computer/runs/computer/results/magic/computer.gds
string GDS_END 88398268
string GDS_START 859364
<< end >>

