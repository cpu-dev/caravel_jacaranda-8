magic
tech sky130A
magscale 1 2
timestamp 1636421769
<< obsli1 >>
rect 1104 2159 390816 391697
<< obsm1 >>
rect 382 1436 391630 391728
<< metal2 >>
rect 1674 393319 1730 394119
rect 5078 393319 5134 394119
rect 8482 393319 8538 394119
rect 11978 393319 12034 394119
rect 15382 393319 15438 394119
rect 18786 393319 18842 394119
rect 22282 393319 22338 394119
rect 25686 393319 25742 394119
rect 29182 393319 29238 394119
rect 32586 393319 32642 394119
rect 35990 393319 36046 394119
rect 39486 393319 39542 394119
rect 42890 393319 42946 394119
rect 46294 393319 46350 394119
rect 49790 393319 49846 394119
rect 53194 393319 53250 394119
rect 56690 393319 56746 394119
rect 60094 393319 60150 394119
rect 63498 393319 63554 394119
rect 66994 393319 67050 394119
rect 70398 393319 70454 394119
rect 73802 393319 73858 394119
rect 77298 393319 77354 394119
rect 80702 393319 80758 394119
rect 84198 393319 84254 394119
rect 87602 393319 87658 394119
rect 91006 393319 91062 394119
rect 94502 393319 94558 394119
rect 97906 393319 97962 394119
rect 101310 393319 101366 394119
rect 104806 393319 104862 394119
rect 108210 393319 108266 394119
rect 111706 393319 111762 394119
rect 115110 393319 115166 394119
rect 118514 393319 118570 394119
rect 122010 393319 122066 394119
rect 125414 393319 125470 394119
rect 128818 393319 128874 394119
rect 132314 393319 132370 394119
rect 135718 393319 135774 394119
rect 139214 393319 139270 394119
rect 142618 393319 142674 394119
rect 146022 393319 146078 394119
rect 149518 393319 149574 394119
rect 152922 393319 152978 394119
rect 156326 393319 156382 394119
rect 159822 393319 159878 394119
rect 163226 393319 163282 394119
rect 166722 393319 166778 394119
rect 170126 393319 170182 394119
rect 173530 393319 173586 394119
rect 177026 393319 177082 394119
rect 180430 393319 180486 394119
rect 183834 393319 183890 394119
rect 187330 393319 187386 394119
rect 190734 393319 190790 394119
rect 194230 393319 194286 394119
rect 197634 393319 197690 394119
rect 201038 393319 201094 394119
rect 204534 393319 204590 394119
rect 207938 393319 207994 394119
rect 211434 393319 211490 394119
rect 214838 393319 214894 394119
rect 218242 393319 218298 394119
rect 221738 393319 221794 394119
rect 225142 393319 225198 394119
rect 228546 393319 228602 394119
rect 232042 393319 232098 394119
rect 235446 393319 235502 394119
rect 238942 393319 238998 394119
rect 242346 393319 242402 394119
rect 245750 393319 245806 394119
rect 249246 393319 249302 394119
rect 252650 393319 252706 394119
rect 256054 393319 256110 394119
rect 259550 393319 259606 394119
rect 262954 393319 263010 394119
rect 266450 393319 266506 394119
rect 269854 393319 269910 394119
rect 273258 393319 273314 394119
rect 276754 393319 276810 394119
rect 280158 393319 280214 394119
rect 283562 393319 283618 394119
rect 287058 393319 287114 394119
rect 290462 393319 290518 394119
rect 293958 393319 294014 394119
rect 297362 393319 297418 394119
rect 300766 393319 300822 394119
rect 304262 393319 304318 394119
rect 307666 393319 307722 394119
rect 311070 393319 311126 394119
rect 314566 393319 314622 394119
rect 317970 393319 318026 394119
rect 321466 393319 321522 394119
rect 324870 393319 324926 394119
rect 328274 393319 328330 394119
rect 331770 393319 331826 394119
rect 335174 393319 335230 394119
rect 338578 393319 338634 394119
rect 342074 393319 342130 394119
rect 345478 393319 345534 394119
rect 348974 393319 349030 394119
rect 352378 393319 352434 394119
rect 355782 393319 355838 394119
rect 359278 393319 359334 394119
rect 362682 393319 362738 394119
rect 366086 393319 366142 394119
rect 369582 393319 369638 394119
rect 372986 393319 373042 394119
rect 376482 393319 376538 394119
rect 379886 393319 379942 394119
rect 383290 393319 383346 394119
rect 386786 393319 386842 394119
rect 390190 393319 390246 394119
rect 386 0 442 800
rect 1122 0 1178 800
rect 1950 0 2006 800
rect 2686 0 2742 800
rect 3514 0 3570 800
rect 4342 0 4398 800
rect 5078 0 5134 800
rect 5906 0 5962 800
rect 6734 0 6790 800
rect 7470 0 7526 800
rect 8298 0 8354 800
rect 9126 0 9182 800
rect 9862 0 9918 800
rect 10690 0 10746 800
rect 11518 0 11574 800
rect 12254 0 12310 800
rect 13082 0 13138 800
rect 13818 0 13874 800
rect 14646 0 14702 800
rect 15474 0 15530 800
rect 16210 0 16266 800
rect 17038 0 17094 800
rect 17866 0 17922 800
rect 18602 0 18658 800
rect 19430 0 19486 800
rect 20258 0 20314 800
rect 20994 0 21050 800
rect 21822 0 21878 800
rect 22650 0 22706 800
rect 23386 0 23442 800
rect 24214 0 24270 800
rect 24950 0 25006 800
rect 25778 0 25834 800
rect 26606 0 26662 800
rect 27342 0 27398 800
rect 28170 0 28226 800
rect 28998 0 29054 800
rect 29734 0 29790 800
rect 30562 0 30618 800
rect 31390 0 31446 800
rect 32126 0 32182 800
rect 32954 0 33010 800
rect 33782 0 33838 800
rect 34518 0 34574 800
rect 35346 0 35402 800
rect 36082 0 36138 800
rect 36910 0 36966 800
rect 37738 0 37794 800
rect 38474 0 38530 800
rect 39302 0 39358 800
rect 40130 0 40186 800
rect 40866 0 40922 800
rect 41694 0 41750 800
rect 42522 0 42578 800
rect 43258 0 43314 800
rect 44086 0 44142 800
rect 44914 0 44970 800
rect 45650 0 45706 800
rect 46478 0 46534 800
rect 47214 0 47270 800
rect 48042 0 48098 800
rect 48870 0 48926 800
rect 49606 0 49662 800
rect 50434 0 50490 800
rect 51262 0 51318 800
rect 51998 0 52054 800
rect 52826 0 52882 800
rect 53654 0 53710 800
rect 54390 0 54446 800
rect 55218 0 55274 800
rect 56046 0 56102 800
rect 56782 0 56838 800
rect 57610 0 57666 800
rect 58346 0 58402 800
rect 59174 0 59230 800
rect 60002 0 60058 800
rect 60738 0 60794 800
rect 61566 0 61622 800
rect 62394 0 62450 800
rect 63130 0 63186 800
rect 63958 0 64014 800
rect 64786 0 64842 800
rect 65522 0 65578 800
rect 66350 0 66406 800
rect 67178 0 67234 800
rect 67914 0 67970 800
rect 68742 0 68798 800
rect 69478 0 69534 800
rect 70306 0 70362 800
rect 71134 0 71190 800
rect 71870 0 71926 800
rect 72698 0 72754 800
rect 73526 0 73582 800
rect 74262 0 74318 800
rect 75090 0 75146 800
rect 75918 0 75974 800
rect 76654 0 76710 800
rect 77482 0 77538 800
rect 78310 0 78366 800
rect 79046 0 79102 800
rect 79874 0 79930 800
rect 80610 0 80666 800
rect 81438 0 81494 800
rect 82266 0 82322 800
rect 83002 0 83058 800
rect 83830 0 83886 800
rect 84658 0 84714 800
rect 85394 0 85450 800
rect 86222 0 86278 800
rect 87050 0 87106 800
rect 87786 0 87842 800
rect 88614 0 88670 800
rect 89442 0 89498 800
rect 90178 0 90234 800
rect 91006 0 91062 800
rect 91742 0 91798 800
rect 92570 0 92626 800
rect 93398 0 93454 800
rect 94134 0 94190 800
rect 94962 0 95018 800
rect 95790 0 95846 800
rect 96526 0 96582 800
rect 97354 0 97410 800
rect 98182 0 98238 800
rect 98918 0 98974 800
rect 99746 0 99802 800
rect 100574 0 100630 800
rect 101310 0 101366 800
rect 102138 0 102194 800
rect 102874 0 102930 800
rect 103702 0 103758 800
rect 104530 0 104586 800
rect 105266 0 105322 800
rect 106094 0 106150 800
rect 106922 0 106978 800
rect 107658 0 107714 800
rect 108486 0 108542 800
rect 109314 0 109370 800
rect 110050 0 110106 800
rect 110878 0 110934 800
rect 111706 0 111762 800
rect 112442 0 112498 800
rect 113270 0 113326 800
rect 114006 0 114062 800
rect 114834 0 114890 800
rect 115662 0 115718 800
rect 116398 0 116454 800
rect 117226 0 117282 800
rect 118054 0 118110 800
rect 118790 0 118846 800
rect 119618 0 119674 800
rect 120446 0 120502 800
rect 121182 0 121238 800
rect 122010 0 122066 800
rect 122838 0 122894 800
rect 123574 0 123630 800
rect 124402 0 124458 800
rect 125138 0 125194 800
rect 125966 0 126022 800
rect 126794 0 126850 800
rect 127530 0 127586 800
rect 128358 0 128414 800
rect 129186 0 129242 800
rect 129922 0 129978 800
rect 130750 0 130806 800
rect 131578 0 131634 800
rect 132314 0 132370 800
rect 133142 0 133198 800
rect 133970 0 134026 800
rect 134706 0 134762 800
rect 135534 0 135590 800
rect 136270 0 136326 800
rect 137098 0 137154 800
rect 137926 0 137982 800
rect 138662 0 138718 800
rect 139490 0 139546 800
rect 140318 0 140374 800
rect 141054 0 141110 800
rect 141882 0 141938 800
rect 142710 0 142766 800
rect 143446 0 143502 800
rect 144274 0 144330 800
rect 145102 0 145158 800
rect 145838 0 145894 800
rect 146666 0 146722 800
rect 147402 0 147458 800
rect 148230 0 148286 800
rect 149058 0 149114 800
rect 149794 0 149850 800
rect 150622 0 150678 800
rect 151450 0 151506 800
rect 152186 0 152242 800
rect 153014 0 153070 800
rect 153842 0 153898 800
rect 154578 0 154634 800
rect 155406 0 155462 800
rect 156234 0 156290 800
rect 156970 0 157026 800
rect 157798 0 157854 800
rect 158534 0 158590 800
rect 159362 0 159418 800
rect 160190 0 160246 800
rect 160926 0 160982 800
rect 161754 0 161810 800
rect 162582 0 162638 800
rect 163318 0 163374 800
rect 164146 0 164202 800
rect 164974 0 165030 800
rect 165710 0 165766 800
rect 166538 0 166594 800
rect 167366 0 167422 800
rect 168102 0 168158 800
rect 168930 0 168986 800
rect 169666 0 169722 800
rect 170494 0 170550 800
rect 171322 0 171378 800
rect 172058 0 172114 800
rect 172886 0 172942 800
rect 173714 0 173770 800
rect 174450 0 174506 800
rect 175278 0 175334 800
rect 176106 0 176162 800
rect 176842 0 176898 800
rect 177670 0 177726 800
rect 178498 0 178554 800
rect 179234 0 179290 800
rect 180062 0 180118 800
rect 180798 0 180854 800
rect 181626 0 181682 800
rect 182454 0 182510 800
rect 183190 0 183246 800
rect 184018 0 184074 800
rect 184846 0 184902 800
rect 185582 0 185638 800
rect 186410 0 186466 800
rect 187238 0 187294 800
rect 187974 0 188030 800
rect 188802 0 188858 800
rect 189630 0 189686 800
rect 190366 0 190422 800
rect 191194 0 191250 800
rect 191930 0 191986 800
rect 192758 0 192814 800
rect 193586 0 193642 800
rect 194322 0 194378 800
rect 195150 0 195206 800
rect 195978 0 196034 800
rect 196714 0 196770 800
rect 197542 0 197598 800
rect 198370 0 198426 800
rect 199106 0 199162 800
rect 199934 0 199990 800
rect 200762 0 200818 800
rect 201498 0 201554 800
rect 202326 0 202382 800
rect 203062 0 203118 800
rect 203890 0 203946 800
rect 204718 0 204774 800
rect 205454 0 205510 800
rect 206282 0 206338 800
rect 207110 0 207166 800
rect 207846 0 207902 800
rect 208674 0 208730 800
rect 209502 0 209558 800
rect 210238 0 210294 800
rect 211066 0 211122 800
rect 211894 0 211950 800
rect 212630 0 212686 800
rect 213458 0 213514 800
rect 214194 0 214250 800
rect 215022 0 215078 800
rect 215850 0 215906 800
rect 216586 0 216642 800
rect 217414 0 217470 800
rect 218242 0 218298 800
rect 218978 0 219034 800
rect 219806 0 219862 800
rect 220634 0 220690 800
rect 221370 0 221426 800
rect 222198 0 222254 800
rect 223026 0 223082 800
rect 223762 0 223818 800
rect 224590 0 224646 800
rect 225326 0 225382 800
rect 226154 0 226210 800
rect 226982 0 227038 800
rect 227718 0 227774 800
rect 228546 0 228602 800
rect 229374 0 229430 800
rect 230110 0 230166 800
rect 230938 0 230994 800
rect 231766 0 231822 800
rect 232502 0 232558 800
rect 233330 0 233386 800
rect 234158 0 234214 800
rect 234894 0 234950 800
rect 235722 0 235778 800
rect 236458 0 236514 800
rect 237286 0 237342 800
rect 238114 0 238170 800
rect 238850 0 238906 800
rect 239678 0 239734 800
rect 240506 0 240562 800
rect 241242 0 241298 800
rect 242070 0 242126 800
rect 242898 0 242954 800
rect 243634 0 243690 800
rect 244462 0 244518 800
rect 245290 0 245346 800
rect 246026 0 246082 800
rect 246854 0 246910 800
rect 247590 0 247646 800
rect 248418 0 248474 800
rect 249246 0 249302 800
rect 249982 0 250038 800
rect 250810 0 250866 800
rect 251638 0 251694 800
rect 252374 0 252430 800
rect 253202 0 253258 800
rect 254030 0 254086 800
rect 254766 0 254822 800
rect 255594 0 255650 800
rect 256422 0 256478 800
rect 257158 0 257214 800
rect 257986 0 258042 800
rect 258722 0 258778 800
rect 259550 0 259606 800
rect 260378 0 260434 800
rect 261114 0 261170 800
rect 261942 0 261998 800
rect 262770 0 262826 800
rect 263506 0 263562 800
rect 264334 0 264390 800
rect 265162 0 265218 800
rect 265898 0 265954 800
rect 266726 0 266782 800
rect 267554 0 267610 800
rect 268290 0 268346 800
rect 269118 0 269174 800
rect 269854 0 269910 800
rect 270682 0 270738 800
rect 271510 0 271566 800
rect 272246 0 272302 800
rect 273074 0 273130 800
rect 273902 0 273958 800
rect 274638 0 274694 800
rect 275466 0 275522 800
rect 276294 0 276350 800
rect 277030 0 277086 800
rect 277858 0 277914 800
rect 278686 0 278742 800
rect 279422 0 279478 800
rect 280250 0 280306 800
rect 280986 0 281042 800
rect 281814 0 281870 800
rect 282642 0 282698 800
rect 283378 0 283434 800
rect 284206 0 284262 800
rect 285034 0 285090 800
rect 285770 0 285826 800
rect 286598 0 286654 800
rect 287426 0 287482 800
rect 288162 0 288218 800
rect 288990 0 289046 800
rect 289818 0 289874 800
rect 290554 0 290610 800
rect 291382 0 291438 800
rect 292118 0 292174 800
rect 292946 0 293002 800
rect 293774 0 293830 800
rect 294510 0 294566 800
rect 295338 0 295394 800
rect 296166 0 296222 800
rect 296902 0 296958 800
rect 297730 0 297786 800
rect 298558 0 298614 800
rect 299294 0 299350 800
rect 300122 0 300178 800
rect 300950 0 301006 800
rect 301686 0 301742 800
rect 302514 0 302570 800
rect 303250 0 303306 800
rect 304078 0 304134 800
rect 304906 0 304962 800
rect 305642 0 305698 800
rect 306470 0 306526 800
rect 307298 0 307354 800
rect 308034 0 308090 800
rect 308862 0 308918 800
rect 309690 0 309746 800
rect 310426 0 310482 800
rect 311254 0 311310 800
rect 312082 0 312138 800
rect 312818 0 312874 800
rect 313646 0 313702 800
rect 314382 0 314438 800
rect 315210 0 315266 800
rect 316038 0 316094 800
rect 316774 0 316830 800
rect 317602 0 317658 800
rect 318430 0 318486 800
rect 319166 0 319222 800
rect 319994 0 320050 800
rect 320822 0 320878 800
rect 321558 0 321614 800
rect 322386 0 322442 800
rect 323214 0 323270 800
rect 323950 0 324006 800
rect 324778 0 324834 800
rect 325514 0 325570 800
rect 326342 0 326398 800
rect 327170 0 327226 800
rect 327906 0 327962 800
rect 328734 0 328790 800
rect 329562 0 329618 800
rect 330298 0 330354 800
rect 331126 0 331182 800
rect 331954 0 332010 800
rect 332690 0 332746 800
rect 333518 0 333574 800
rect 334346 0 334402 800
rect 335082 0 335138 800
rect 335910 0 335966 800
rect 336646 0 336702 800
rect 337474 0 337530 800
rect 338302 0 338358 800
rect 339038 0 339094 800
rect 339866 0 339922 800
rect 340694 0 340750 800
rect 341430 0 341486 800
rect 342258 0 342314 800
rect 343086 0 343142 800
rect 343822 0 343878 800
rect 344650 0 344706 800
rect 345478 0 345534 800
rect 346214 0 346270 800
rect 347042 0 347098 800
rect 347778 0 347834 800
rect 348606 0 348662 800
rect 349434 0 349490 800
rect 350170 0 350226 800
rect 350998 0 351054 800
rect 351826 0 351882 800
rect 352562 0 352618 800
rect 353390 0 353446 800
rect 354218 0 354274 800
rect 354954 0 355010 800
rect 355782 0 355838 800
rect 356610 0 356666 800
rect 357346 0 357402 800
rect 358174 0 358230 800
rect 358910 0 358966 800
rect 359738 0 359794 800
rect 360566 0 360622 800
rect 361302 0 361358 800
rect 362130 0 362186 800
rect 362958 0 363014 800
rect 363694 0 363750 800
rect 364522 0 364578 800
rect 365350 0 365406 800
rect 366086 0 366142 800
rect 366914 0 366970 800
rect 367742 0 367798 800
rect 368478 0 368534 800
rect 369306 0 369362 800
rect 370042 0 370098 800
rect 370870 0 370926 800
rect 371698 0 371754 800
rect 372434 0 372490 800
rect 373262 0 373318 800
rect 374090 0 374146 800
rect 374826 0 374882 800
rect 375654 0 375710 800
rect 376482 0 376538 800
rect 377218 0 377274 800
rect 378046 0 378102 800
rect 378874 0 378930 800
rect 379610 0 379666 800
rect 380438 0 380494 800
rect 381174 0 381230 800
rect 382002 0 382058 800
rect 382830 0 382886 800
rect 383566 0 383622 800
rect 384394 0 384450 800
rect 385222 0 385278 800
rect 385958 0 386014 800
rect 386786 0 386842 800
rect 387614 0 387670 800
rect 388350 0 388406 800
rect 389178 0 389234 800
rect 390006 0 390062 800
rect 390742 0 390798 800
rect 391570 0 391626 800
<< obsm2 >>
rect 388 393263 1618 393319
rect 1786 393263 5022 393319
rect 5190 393263 8426 393319
rect 8594 393263 11922 393319
rect 12090 393263 15326 393319
rect 15494 393263 18730 393319
rect 18898 393263 22226 393319
rect 22394 393263 25630 393319
rect 25798 393263 29126 393319
rect 29294 393263 32530 393319
rect 32698 393263 35934 393319
rect 36102 393263 39430 393319
rect 39598 393263 42834 393319
rect 43002 393263 46238 393319
rect 46406 393263 49734 393319
rect 49902 393263 53138 393319
rect 53306 393263 56634 393319
rect 56802 393263 60038 393319
rect 60206 393263 63442 393319
rect 63610 393263 66938 393319
rect 67106 393263 70342 393319
rect 70510 393263 73746 393319
rect 73914 393263 77242 393319
rect 77410 393263 80646 393319
rect 80814 393263 84142 393319
rect 84310 393263 87546 393319
rect 87714 393263 90950 393319
rect 91118 393263 94446 393319
rect 94614 393263 97850 393319
rect 98018 393263 101254 393319
rect 101422 393263 104750 393319
rect 104918 393263 108154 393319
rect 108322 393263 111650 393319
rect 111818 393263 115054 393319
rect 115222 393263 118458 393319
rect 118626 393263 121954 393319
rect 122122 393263 125358 393319
rect 125526 393263 128762 393319
rect 128930 393263 132258 393319
rect 132426 393263 135662 393319
rect 135830 393263 139158 393319
rect 139326 393263 142562 393319
rect 142730 393263 145966 393319
rect 146134 393263 149462 393319
rect 149630 393263 152866 393319
rect 153034 393263 156270 393319
rect 156438 393263 159766 393319
rect 159934 393263 163170 393319
rect 163338 393263 166666 393319
rect 166834 393263 170070 393319
rect 170238 393263 173474 393319
rect 173642 393263 176970 393319
rect 177138 393263 180374 393319
rect 180542 393263 183778 393319
rect 183946 393263 187274 393319
rect 187442 393263 190678 393319
rect 190846 393263 194174 393319
rect 194342 393263 197578 393319
rect 197746 393263 200982 393319
rect 201150 393263 204478 393319
rect 204646 393263 207882 393319
rect 208050 393263 211378 393319
rect 211546 393263 214782 393319
rect 214950 393263 218186 393319
rect 218354 393263 221682 393319
rect 221850 393263 225086 393319
rect 225254 393263 228490 393319
rect 228658 393263 231986 393319
rect 232154 393263 235390 393319
rect 235558 393263 238886 393319
rect 239054 393263 242290 393319
rect 242458 393263 245694 393319
rect 245862 393263 249190 393319
rect 249358 393263 252594 393319
rect 252762 393263 255998 393319
rect 256166 393263 259494 393319
rect 259662 393263 262898 393319
rect 263066 393263 266394 393319
rect 266562 393263 269798 393319
rect 269966 393263 273202 393319
rect 273370 393263 276698 393319
rect 276866 393263 280102 393319
rect 280270 393263 283506 393319
rect 283674 393263 287002 393319
rect 287170 393263 290406 393319
rect 290574 393263 293902 393319
rect 294070 393263 297306 393319
rect 297474 393263 300710 393319
rect 300878 393263 304206 393319
rect 304374 393263 307610 393319
rect 307778 393263 311014 393319
rect 311182 393263 314510 393319
rect 314678 393263 317914 393319
rect 318082 393263 321410 393319
rect 321578 393263 324814 393319
rect 324982 393263 328218 393319
rect 328386 393263 331714 393319
rect 331882 393263 335118 393319
rect 335286 393263 338522 393319
rect 338690 393263 342018 393319
rect 342186 393263 345422 393319
rect 345590 393263 348918 393319
rect 349086 393263 352322 393319
rect 352490 393263 355726 393319
rect 355894 393263 359222 393319
rect 359390 393263 362626 393319
rect 362794 393263 366030 393319
rect 366198 393263 369526 393319
rect 369694 393263 372930 393319
rect 373098 393263 376426 393319
rect 376594 393263 379830 393319
rect 379998 393263 383234 393319
rect 383402 393263 386730 393319
rect 386898 393263 390134 393319
rect 390302 393263 391624 393319
rect 388 856 391624 393263
rect 498 734 1066 856
rect 1234 734 1894 856
rect 2062 734 2630 856
rect 2798 734 3458 856
rect 3626 734 4286 856
rect 4454 734 5022 856
rect 5190 734 5850 856
rect 6018 734 6678 856
rect 6846 734 7414 856
rect 7582 734 8242 856
rect 8410 734 9070 856
rect 9238 734 9806 856
rect 9974 734 10634 856
rect 10802 734 11462 856
rect 11630 734 12198 856
rect 12366 734 13026 856
rect 13194 734 13762 856
rect 13930 734 14590 856
rect 14758 734 15418 856
rect 15586 734 16154 856
rect 16322 734 16982 856
rect 17150 734 17810 856
rect 17978 734 18546 856
rect 18714 734 19374 856
rect 19542 734 20202 856
rect 20370 734 20938 856
rect 21106 734 21766 856
rect 21934 734 22594 856
rect 22762 734 23330 856
rect 23498 734 24158 856
rect 24326 734 24894 856
rect 25062 734 25722 856
rect 25890 734 26550 856
rect 26718 734 27286 856
rect 27454 734 28114 856
rect 28282 734 28942 856
rect 29110 734 29678 856
rect 29846 734 30506 856
rect 30674 734 31334 856
rect 31502 734 32070 856
rect 32238 734 32898 856
rect 33066 734 33726 856
rect 33894 734 34462 856
rect 34630 734 35290 856
rect 35458 734 36026 856
rect 36194 734 36854 856
rect 37022 734 37682 856
rect 37850 734 38418 856
rect 38586 734 39246 856
rect 39414 734 40074 856
rect 40242 734 40810 856
rect 40978 734 41638 856
rect 41806 734 42466 856
rect 42634 734 43202 856
rect 43370 734 44030 856
rect 44198 734 44858 856
rect 45026 734 45594 856
rect 45762 734 46422 856
rect 46590 734 47158 856
rect 47326 734 47986 856
rect 48154 734 48814 856
rect 48982 734 49550 856
rect 49718 734 50378 856
rect 50546 734 51206 856
rect 51374 734 51942 856
rect 52110 734 52770 856
rect 52938 734 53598 856
rect 53766 734 54334 856
rect 54502 734 55162 856
rect 55330 734 55990 856
rect 56158 734 56726 856
rect 56894 734 57554 856
rect 57722 734 58290 856
rect 58458 734 59118 856
rect 59286 734 59946 856
rect 60114 734 60682 856
rect 60850 734 61510 856
rect 61678 734 62338 856
rect 62506 734 63074 856
rect 63242 734 63902 856
rect 64070 734 64730 856
rect 64898 734 65466 856
rect 65634 734 66294 856
rect 66462 734 67122 856
rect 67290 734 67858 856
rect 68026 734 68686 856
rect 68854 734 69422 856
rect 69590 734 70250 856
rect 70418 734 71078 856
rect 71246 734 71814 856
rect 71982 734 72642 856
rect 72810 734 73470 856
rect 73638 734 74206 856
rect 74374 734 75034 856
rect 75202 734 75862 856
rect 76030 734 76598 856
rect 76766 734 77426 856
rect 77594 734 78254 856
rect 78422 734 78990 856
rect 79158 734 79818 856
rect 79986 734 80554 856
rect 80722 734 81382 856
rect 81550 734 82210 856
rect 82378 734 82946 856
rect 83114 734 83774 856
rect 83942 734 84602 856
rect 84770 734 85338 856
rect 85506 734 86166 856
rect 86334 734 86994 856
rect 87162 734 87730 856
rect 87898 734 88558 856
rect 88726 734 89386 856
rect 89554 734 90122 856
rect 90290 734 90950 856
rect 91118 734 91686 856
rect 91854 734 92514 856
rect 92682 734 93342 856
rect 93510 734 94078 856
rect 94246 734 94906 856
rect 95074 734 95734 856
rect 95902 734 96470 856
rect 96638 734 97298 856
rect 97466 734 98126 856
rect 98294 734 98862 856
rect 99030 734 99690 856
rect 99858 734 100518 856
rect 100686 734 101254 856
rect 101422 734 102082 856
rect 102250 734 102818 856
rect 102986 734 103646 856
rect 103814 734 104474 856
rect 104642 734 105210 856
rect 105378 734 106038 856
rect 106206 734 106866 856
rect 107034 734 107602 856
rect 107770 734 108430 856
rect 108598 734 109258 856
rect 109426 734 109994 856
rect 110162 734 110822 856
rect 110990 734 111650 856
rect 111818 734 112386 856
rect 112554 734 113214 856
rect 113382 734 113950 856
rect 114118 734 114778 856
rect 114946 734 115606 856
rect 115774 734 116342 856
rect 116510 734 117170 856
rect 117338 734 117998 856
rect 118166 734 118734 856
rect 118902 734 119562 856
rect 119730 734 120390 856
rect 120558 734 121126 856
rect 121294 734 121954 856
rect 122122 734 122782 856
rect 122950 734 123518 856
rect 123686 734 124346 856
rect 124514 734 125082 856
rect 125250 734 125910 856
rect 126078 734 126738 856
rect 126906 734 127474 856
rect 127642 734 128302 856
rect 128470 734 129130 856
rect 129298 734 129866 856
rect 130034 734 130694 856
rect 130862 734 131522 856
rect 131690 734 132258 856
rect 132426 734 133086 856
rect 133254 734 133914 856
rect 134082 734 134650 856
rect 134818 734 135478 856
rect 135646 734 136214 856
rect 136382 734 137042 856
rect 137210 734 137870 856
rect 138038 734 138606 856
rect 138774 734 139434 856
rect 139602 734 140262 856
rect 140430 734 140998 856
rect 141166 734 141826 856
rect 141994 734 142654 856
rect 142822 734 143390 856
rect 143558 734 144218 856
rect 144386 734 145046 856
rect 145214 734 145782 856
rect 145950 734 146610 856
rect 146778 734 147346 856
rect 147514 734 148174 856
rect 148342 734 149002 856
rect 149170 734 149738 856
rect 149906 734 150566 856
rect 150734 734 151394 856
rect 151562 734 152130 856
rect 152298 734 152958 856
rect 153126 734 153786 856
rect 153954 734 154522 856
rect 154690 734 155350 856
rect 155518 734 156178 856
rect 156346 734 156914 856
rect 157082 734 157742 856
rect 157910 734 158478 856
rect 158646 734 159306 856
rect 159474 734 160134 856
rect 160302 734 160870 856
rect 161038 734 161698 856
rect 161866 734 162526 856
rect 162694 734 163262 856
rect 163430 734 164090 856
rect 164258 734 164918 856
rect 165086 734 165654 856
rect 165822 734 166482 856
rect 166650 734 167310 856
rect 167478 734 168046 856
rect 168214 734 168874 856
rect 169042 734 169610 856
rect 169778 734 170438 856
rect 170606 734 171266 856
rect 171434 734 172002 856
rect 172170 734 172830 856
rect 172998 734 173658 856
rect 173826 734 174394 856
rect 174562 734 175222 856
rect 175390 734 176050 856
rect 176218 734 176786 856
rect 176954 734 177614 856
rect 177782 734 178442 856
rect 178610 734 179178 856
rect 179346 734 180006 856
rect 180174 734 180742 856
rect 180910 734 181570 856
rect 181738 734 182398 856
rect 182566 734 183134 856
rect 183302 734 183962 856
rect 184130 734 184790 856
rect 184958 734 185526 856
rect 185694 734 186354 856
rect 186522 734 187182 856
rect 187350 734 187918 856
rect 188086 734 188746 856
rect 188914 734 189574 856
rect 189742 734 190310 856
rect 190478 734 191138 856
rect 191306 734 191874 856
rect 192042 734 192702 856
rect 192870 734 193530 856
rect 193698 734 194266 856
rect 194434 734 195094 856
rect 195262 734 195922 856
rect 196090 734 196658 856
rect 196826 734 197486 856
rect 197654 734 198314 856
rect 198482 734 199050 856
rect 199218 734 199878 856
rect 200046 734 200706 856
rect 200874 734 201442 856
rect 201610 734 202270 856
rect 202438 734 203006 856
rect 203174 734 203834 856
rect 204002 734 204662 856
rect 204830 734 205398 856
rect 205566 734 206226 856
rect 206394 734 207054 856
rect 207222 734 207790 856
rect 207958 734 208618 856
rect 208786 734 209446 856
rect 209614 734 210182 856
rect 210350 734 211010 856
rect 211178 734 211838 856
rect 212006 734 212574 856
rect 212742 734 213402 856
rect 213570 734 214138 856
rect 214306 734 214966 856
rect 215134 734 215794 856
rect 215962 734 216530 856
rect 216698 734 217358 856
rect 217526 734 218186 856
rect 218354 734 218922 856
rect 219090 734 219750 856
rect 219918 734 220578 856
rect 220746 734 221314 856
rect 221482 734 222142 856
rect 222310 734 222970 856
rect 223138 734 223706 856
rect 223874 734 224534 856
rect 224702 734 225270 856
rect 225438 734 226098 856
rect 226266 734 226926 856
rect 227094 734 227662 856
rect 227830 734 228490 856
rect 228658 734 229318 856
rect 229486 734 230054 856
rect 230222 734 230882 856
rect 231050 734 231710 856
rect 231878 734 232446 856
rect 232614 734 233274 856
rect 233442 734 234102 856
rect 234270 734 234838 856
rect 235006 734 235666 856
rect 235834 734 236402 856
rect 236570 734 237230 856
rect 237398 734 238058 856
rect 238226 734 238794 856
rect 238962 734 239622 856
rect 239790 734 240450 856
rect 240618 734 241186 856
rect 241354 734 242014 856
rect 242182 734 242842 856
rect 243010 734 243578 856
rect 243746 734 244406 856
rect 244574 734 245234 856
rect 245402 734 245970 856
rect 246138 734 246798 856
rect 246966 734 247534 856
rect 247702 734 248362 856
rect 248530 734 249190 856
rect 249358 734 249926 856
rect 250094 734 250754 856
rect 250922 734 251582 856
rect 251750 734 252318 856
rect 252486 734 253146 856
rect 253314 734 253974 856
rect 254142 734 254710 856
rect 254878 734 255538 856
rect 255706 734 256366 856
rect 256534 734 257102 856
rect 257270 734 257930 856
rect 258098 734 258666 856
rect 258834 734 259494 856
rect 259662 734 260322 856
rect 260490 734 261058 856
rect 261226 734 261886 856
rect 262054 734 262714 856
rect 262882 734 263450 856
rect 263618 734 264278 856
rect 264446 734 265106 856
rect 265274 734 265842 856
rect 266010 734 266670 856
rect 266838 734 267498 856
rect 267666 734 268234 856
rect 268402 734 269062 856
rect 269230 734 269798 856
rect 269966 734 270626 856
rect 270794 734 271454 856
rect 271622 734 272190 856
rect 272358 734 273018 856
rect 273186 734 273846 856
rect 274014 734 274582 856
rect 274750 734 275410 856
rect 275578 734 276238 856
rect 276406 734 276974 856
rect 277142 734 277802 856
rect 277970 734 278630 856
rect 278798 734 279366 856
rect 279534 734 280194 856
rect 280362 734 280930 856
rect 281098 734 281758 856
rect 281926 734 282586 856
rect 282754 734 283322 856
rect 283490 734 284150 856
rect 284318 734 284978 856
rect 285146 734 285714 856
rect 285882 734 286542 856
rect 286710 734 287370 856
rect 287538 734 288106 856
rect 288274 734 288934 856
rect 289102 734 289762 856
rect 289930 734 290498 856
rect 290666 734 291326 856
rect 291494 734 292062 856
rect 292230 734 292890 856
rect 293058 734 293718 856
rect 293886 734 294454 856
rect 294622 734 295282 856
rect 295450 734 296110 856
rect 296278 734 296846 856
rect 297014 734 297674 856
rect 297842 734 298502 856
rect 298670 734 299238 856
rect 299406 734 300066 856
rect 300234 734 300894 856
rect 301062 734 301630 856
rect 301798 734 302458 856
rect 302626 734 303194 856
rect 303362 734 304022 856
rect 304190 734 304850 856
rect 305018 734 305586 856
rect 305754 734 306414 856
rect 306582 734 307242 856
rect 307410 734 307978 856
rect 308146 734 308806 856
rect 308974 734 309634 856
rect 309802 734 310370 856
rect 310538 734 311198 856
rect 311366 734 312026 856
rect 312194 734 312762 856
rect 312930 734 313590 856
rect 313758 734 314326 856
rect 314494 734 315154 856
rect 315322 734 315982 856
rect 316150 734 316718 856
rect 316886 734 317546 856
rect 317714 734 318374 856
rect 318542 734 319110 856
rect 319278 734 319938 856
rect 320106 734 320766 856
rect 320934 734 321502 856
rect 321670 734 322330 856
rect 322498 734 323158 856
rect 323326 734 323894 856
rect 324062 734 324722 856
rect 324890 734 325458 856
rect 325626 734 326286 856
rect 326454 734 327114 856
rect 327282 734 327850 856
rect 328018 734 328678 856
rect 328846 734 329506 856
rect 329674 734 330242 856
rect 330410 734 331070 856
rect 331238 734 331898 856
rect 332066 734 332634 856
rect 332802 734 333462 856
rect 333630 734 334290 856
rect 334458 734 335026 856
rect 335194 734 335854 856
rect 336022 734 336590 856
rect 336758 734 337418 856
rect 337586 734 338246 856
rect 338414 734 338982 856
rect 339150 734 339810 856
rect 339978 734 340638 856
rect 340806 734 341374 856
rect 341542 734 342202 856
rect 342370 734 343030 856
rect 343198 734 343766 856
rect 343934 734 344594 856
rect 344762 734 345422 856
rect 345590 734 346158 856
rect 346326 734 346986 856
rect 347154 734 347722 856
rect 347890 734 348550 856
rect 348718 734 349378 856
rect 349546 734 350114 856
rect 350282 734 350942 856
rect 351110 734 351770 856
rect 351938 734 352506 856
rect 352674 734 353334 856
rect 353502 734 354162 856
rect 354330 734 354898 856
rect 355066 734 355726 856
rect 355894 734 356554 856
rect 356722 734 357290 856
rect 357458 734 358118 856
rect 358286 734 358854 856
rect 359022 734 359682 856
rect 359850 734 360510 856
rect 360678 734 361246 856
rect 361414 734 362074 856
rect 362242 734 362902 856
rect 363070 734 363638 856
rect 363806 734 364466 856
rect 364634 734 365294 856
rect 365462 734 366030 856
rect 366198 734 366858 856
rect 367026 734 367686 856
rect 367854 734 368422 856
rect 368590 734 369250 856
rect 369418 734 369986 856
rect 370154 734 370814 856
rect 370982 734 371642 856
rect 371810 734 372378 856
rect 372546 734 373206 856
rect 373374 734 374034 856
rect 374202 734 374770 856
rect 374938 734 375598 856
rect 375766 734 376426 856
rect 376594 734 377162 856
rect 377330 734 377990 856
rect 378158 734 378818 856
rect 378986 734 379554 856
rect 379722 734 380382 856
rect 380550 734 381118 856
rect 381286 734 381946 856
rect 382114 734 382774 856
rect 382942 734 383510 856
rect 383678 734 384338 856
rect 384506 734 385166 856
rect 385334 734 385902 856
rect 386070 734 386730 856
rect 386898 734 387558 856
rect 387726 734 388294 856
rect 388462 734 389122 856
rect 389290 734 389950 856
rect 390118 734 390686 856
rect 390854 734 391514 856
<< obsm3 >>
rect 4208 2143 388528 391713
<< metal4 >>
rect 4208 2128 4528 391728
rect 19568 2128 19888 391728
rect 34928 2128 35248 391728
rect 50288 2128 50608 391728
rect 65648 2128 65968 391728
rect 81008 2128 81328 391728
rect 96368 2128 96688 391728
rect 111728 2128 112048 391728
rect 127088 2128 127408 391728
rect 142448 2128 142768 391728
rect 157808 2128 158128 391728
rect 173168 2128 173488 391728
rect 188528 2128 188848 391728
rect 203888 2128 204208 391728
rect 219248 2128 219568 391728
rect 234608 2128 234928 391728
rect 249968 2128 250288 391728
rect 265328 2128 265648 391728
rect 280688 2128 281008 391728
rect 296048 2128 296368 391728
rect 311408 2128 311728 391728
rect 326768 2128 327088 391728
rect 342128 2128 342448 391728
rect 357488 2128 357808 391728
rect 372848 2128 373168 391728
rect 388208 2128 388528 391728
<< obsm4 >>
rect 120763 214643 121013 215661
<< labels >>
rlabel metal2 s 1674 393319 1730 394119 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 104806 393319 104862 394119 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 115110 393319 115166 394119 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 125414 393319 125470 394119 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 135718 393319 135774 394119 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 146022 393319 146078 394119 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 156326 393319 156382 394119 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 166722 393319 166778 394119 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 177026 393319 177082 394119 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 187330 393319 187386 394119 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 197634 393319 197690 394119 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 11978 393319 12034 394119 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 207938 393319 207994 394119 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 218242 393319 218298 394119 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 228546 393319 228602 394119 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 238942 393319 238998 394119 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 249246 393319 249302 394119 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 259550 393319 259606 394119 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 269854 393319 269910 394119 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 280158 393319 280214 394119 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 290462 393319 290518 394119 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 300766 393319 300822 394119 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 22282 393319 22338 394119 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 311070 393319 311126 394119 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 321466 393319 321522 394119 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 331770 393319 331826 394119 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 342074 393319 342130 394119 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 352378 393319 352434 394119 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 362682 393319 362738 394119 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 372986 393319 373042 394119 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 383290 393319 383346 394119 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 32586 393319 32642 394119 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 42890 393319 42946 394119 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 53194 393319 53250 394119 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 63498 393319 63554 394119 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 73802 393319 73858 394119 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 84198 393319 84254 394119 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 94502 393319 94558 394119 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5078 393319 5134 394119 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 108210 393319 108266 394119 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 118514 393319 118570 394119 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 128818 393319 128874 394119 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 139214 393319 139270 394119 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 149518 393319 149574 394119 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 159822 393319 159878 394119 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 170126 393319 170182 394119 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 180430 393319 180486 394119 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 190734 393319 190790 394119 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 201038 393319 201094 394119 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 15382 393319 15438 394119 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 211434 393319 211490 394119 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 221738 393319 221794 394119 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 232042 393319 232098 394119 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 242346 393319 242402 394119 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 252650 393319 252706 394119 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 262954 393319 263010 394119 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 273258 393319 273314 394119 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 283562 393319 283618 394119 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 293958 393319 294014 394119 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 304262 393319 304318 394119 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 25686 393319 25742 394119 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 314566 393319 314622 394119 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 324870 393319 324926 394119 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 335174 393319 335230 394119 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 345478 393319 345534 394119 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 355782 393319 355838 394119 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 366086 393319 366142 394119 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 376482 393319 376538 394119 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 386786 393319 386842 394119 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 35990 393319 36046 394119 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 46294 393319 46350 394119 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 56690 393319 56746 394119 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 66994 393319 67050 394119 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 77298 393319 77354 394119 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 87602 393319 87658 394119 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 97906 393319 97962 394119 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 8482 393319 8538 394119 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 111706 393319 111762 394119 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 122010 393319 122066 394119 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 132314 393319 132370 394119 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 142618 393319 142674 394119 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 152922 393319 152978 394119 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 163226 393319 163282 394119 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 173530 393319 173586 394119 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 183834 393319 183890 394119 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 194230 393319 194286 394119 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 204534 393319 204590 394119 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 18786 393319 18842 394119 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 214838 393319 214894 394119 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 225142 393319 225198 394119 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 235446 393319 235502 394119 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 245750 393319 245806 394119 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 256054 393319 256110 394119 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 266450 393319 266506 394119 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 276754 393319 276810 394119 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 287058 393319 287114 394119 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 297362 393319 297418 394119 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 307666 393319 307722 394119 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 29182 393319 29238 394119 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 317970 393319 318026 394119 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 328274 393319 328330 394119 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 338578 393319 338634 394119 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 348974 393319 349030 394119 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 359278 393319 359334 394119 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 369582 393319 369638 394119 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 379886 393319 379942 394119 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 390190 393319 390246 394119 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 39486 393319 39542 394119 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 49790 393319 49846 394119 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 60094 393319 60150 394119 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 70398 393319 70454 394119 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 80702 393319 80758 394119 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 91006 393319 91062 394119 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 101310 393319 101366 394119 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 390006 0 390062 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 390742 0 390798 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 391570 0 391626 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 323214 0 323270 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 325514 0 325570 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 327906 0 327962 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 330298 0 330354 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 332690 0 332746 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 335082 0 335138 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 337474 0 337530 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 339866 0 339922 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 342258 0 342314 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 344650 0 344706 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 347042 0 347098 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 349434 0 349490 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 351826 0 351882 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 354218 0 354274 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 356610 0 356666 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 358910 0 358966 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 361302 0 361358 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 363694 0 363750 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 366086 0 366142 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 368478 0 368534 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 370870 0 370926 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 373262 0 373318 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 375654 0 375710 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 378046 0 378102 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 380438 0 380494 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 382830 0 382886 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 385222 0 385278 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 387614 0 387670 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 170494 0 170550 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 182454 0 182510 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 184846 0 184902 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 194322 0 194378 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 196714 0 196770 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 203890 0 203946 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 206282 0 206338 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 211066 0 211122 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 215850 0 215906 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 220634 0 220690 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 223026 0 223082 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 225326 0 225382 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 227718 0 227774 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 230110 0 230166 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 234894 0 234950 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 237286 0 237342 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 242070 0 242126 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 244462 0 244518 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 246854 0 246910 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 249246 0 249302 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 251638 0 251694 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 254030 0 254086 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 256422 0 256478 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 258722 0 258778 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 261114 0 261170 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 263506 0 263562 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 265898 0 265954 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 268290 0 268346 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 270682 0 270738 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 273074 0 273130 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 275466 0 275522 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 277858 0 277914 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 280250 0 280306 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 282642 0 282698 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 285034 0 285090 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 287426 0 287482 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 289818 0 289874 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 292118 0 292174 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 294510 0 294566 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 296902 0 296958 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 299294 0 299350 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 301686 0 301742 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 304078 0 304134 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 306470 0 306526 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 308862 0 308918 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 311254 0 311310 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 313646 0 313702 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 316038 0 316094 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 318430 0 318486 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 320822 0 320878 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 323950 0 324006 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 326342 0 326398 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 328734 0 328790 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 331126 0 331182 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 333518 0 333574 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 335910 0 335966 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 338302 0 338358 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 340694 0 340750 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 343086 0 343142 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 345478 0 345534 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 347778 0 347834 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 350170 0 350226 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 352562 0 352618 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 354954 0 355010 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 357346 0 357402 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 359738 0 359794 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 362130 0 362186 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 364522 0 364578 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 366914 0 366970 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 369306 0 369362 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 371698 0 371754 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 374090 0 374146 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 376482 0 376538 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 378874 0 378930 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 381174 0 381230 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 383566 0 383622 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 385958 0 386014 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 388350 0 388406 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 128358 0 128414 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 142710 0 142766 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 145102 0 145158 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 149794 0 149850 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 152186 0 152242 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 161754 0 161810 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 164146 0 164202 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 173714 0 173770 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 176106 0 176162 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 178498 0 178554 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 180798 0 180854 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 185582 0 185638 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 187974 0 188030 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 190366 0 190422 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 192758 0 192814 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 195150 0 195206 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 197542 0 197598 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 199934 0 199990 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 202326 0 202382 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 204718 0 204774 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 207110 0 207166 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 209502 0 209558 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 211894 0 211950 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 214194 0 214250 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 216586 0 216642 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 218978 0 219034 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 221370 0 221426 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 223762 0 223818 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 226154 0 226210 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 228546 0 228602 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 230938 0 230994 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 233330 0 233386 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 235722 0 235778 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 238114 0 238170 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 240506 0 240562 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 242898 0 242954 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 245290 0 245346 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 247590 0 247646 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 249982 0 250038 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 99746 0 99802 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 252374 0 252430 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 254766 0 254822 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 257158 0 257214 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 259550 0 259606 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 261942 0 261998 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 264334 0 264390 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 266726 0 266782 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 269118 0 269174 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 271510 0 271566 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 273902 0 273958 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 276294 0 276350 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 278686 0 278742 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 280986 0 281042 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 283378 0 283434 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 285770 0 285826 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 288162 0 288218 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 290554 0 290610 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 292946 0 293002 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 295338 0 295394 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 297730 0 297786 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 300122 0 300178 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 302514 0 302570 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 304906 0 304962 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 307298 0 307354 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 309690 0 309746 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 312082 0 312138 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 314382 0 314438 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 316774 0 316830 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 319166 0 319222 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 321558 0 321614 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 324778 0 324834 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 327170 0 327226 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 329562 0 329618 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 331954 0 332010 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 334346 0 334402 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 336646 0 336702 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 339038 0 339094 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 341430 0 341486 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 343822 0 343878 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 346214 0 346270 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 348606 0 348662 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 350998 0 351054 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 353390 0 353446 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 355782 0 355838 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 358174 0 358230 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 360566 0 360622 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 362958 0 363014 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 365350 0 365406 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 367742 0 367798 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 370042 0 370098 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 372434 0 372490 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 374826 0 374882 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 377218 0 377274 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 379610 0 379666 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 382002 0 382058 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 384394 0 384450 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 386786 0 386842 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 389178 0 389234 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 181626 0 181682 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 184018 0 184074 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 186410 0 186466 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 193586 0 193642 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 198370 0 198426 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 200762 0 200818 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 207846 0 207902 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 210238 0 210294 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 212630 0 212686 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 217414 0 217470 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 219806 0 219862 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 224590 0 224646 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 226982 0 227038 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 229374 0 229430 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 231766 0 231822 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 234158 0 234214 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 236458 0 236514 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 241242 0 241298 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 243634 0 243690 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 248418 0 248474 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 250810 0 250866 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 253202 0 253258 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 255594 0 255650 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 257986 0 258042 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 260378 0 260434 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 262770 0 262826 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 265162 0 265218 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 267554 0 267610 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 269854 0 269910 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 272246 0 272302 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 274638 0 274694 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 277030 0 277086 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 279422 0 279478 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 281814 0 281870 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 284206 0 284262 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 286598 0 286654 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 288990 0 289046 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 291382 0 291438 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 293774 0 293830 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 296166 0 296222 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 298558 0 298614 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 300950 0 301006 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 303250 0 303306 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 305642 0 305698 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 308034 0 308090 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 310426 0 310482 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 312818 0 312874 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 317602 0 317658 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 319994 0 320050 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 322386 0 322442 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 391728 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 391728 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 391728 6 vssd1
port 503 nsew ground input
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 391975 394119
string LEFview TRUE
string GDS_FILE /project/openlane/computer/runs/computer/results/magic/computer.gds
string GDS_END 95035594
string GDS_START 1246144
<< end >>

